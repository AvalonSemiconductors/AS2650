// This is the unpowered netlist.
module wrapped_as2650 (wb_clk_i,
    wb_rst_i,
    io_in,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 input [37:0] io_in;
 output [37:0] io_oeb;
 output [37:0] io_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire \as2650.addr_buff[0] ;
 wire \as2650.addr_buff[1] ;
 wire \as2650.addr_buff[2] ;
 wire \as2650.addr_buff[3] ;
 wire \as2650.addr_buff[4] ;
 wire \as2650.addr_buff[5] ;
 wire \as2650.addr_buff[6] ;
 wire \as2650.addr_buff[7] ;
 wire \as2650.carry ;
 wire \as2650.cycle[0] ;
 wire \as2650.cycle[1] ;
 wire \as2650.cycle[2] ;
 wire \as2650.cycle[3] ;
 wire \as2650.cycle[4] ;
 wire \as2650.cycle[5] ;
 wire \as2650.cycle[6] ;
 wire \as2650.cycle[7] ;
 wire \as2650.halted ;
 wire \as2650.holding_reg[0] ;
 wire \as2650.holding_reg[1] ;
 wire \as2650.holding_reg[2] ;
 wire \as2650.holding_reg[3] ;
 wire \as2650.holding_reg[4] ;
 wire \as2650.holding_reg[5] ;
 wire \as2650.holding_reg[6] ;
 wire \as2650.holding_reg[7] ;
 wire \as2650.idx_ctrl[0] ;
 wire \as2650.idx_ctrl[1] ;
 wire \as2650.ins_reg[0] ;
 wire \as2650.ins_reg[1] ;
 wire \as2650.ins_reg[2] ;
 wire \as2650.ins_reg[3] ;
 wire \as2650.ins_reg[4] ;
 wire \as2650.ins_reg[5] ;
 wire \as2650.ins_reg[6] ;
 wire \as2650.ins_reg[7] ;
 wire \as2650.overflow ;
 wire \as2650.pc[0] ;
 wire \as2650.pc[10] ;
 wire \as2650.pc[11] ;
 wire \as2650.pc[12] ;
 wire \as2650.pc[1] ;
 wire \as2650.pc[2] ;
 wire \as2650.pc[3] ;
 wire \as2650.pc[4] ;
 wire \as2650.pc[5] ;
 wire \as2650.pc[6] ;
 wire \as2650.pc[7] ;
 wire \as2650.pc[8] ;
 wire \as2650.pc[9] ;
 wire \as2650.psl[1] ;
 wire \as2650.psl[3] ;
 wire \as2650.psl[4] ;
 wire \as2650.psl[5] ;
 wire \as2650.psl[6] ;
 wire \as2650.psl[7] ;
 wire \as2650.psu[0] ;
 wire \as2650.psu[1] ;
 wire \as2650.psu[2] ;
 wire \as2650.psu[3] ;
 wire \as2650.psu[4] ;
 wire \as2650.psu[5] ;
 wire \as2650.psu[7] ;
 wire \as2650.r0[0] ;
 wire \as2650.r0[1] ;
 wire \as2650.r0[2] ;
 wire \as2650.r0[3] ;
 wire \as2650.r0[4] ;
 wire \as2650.r0[5] ;
 wire \as2650.r0[6] ;
 wire \as2650.r0[7] ;
 wire \as2650.r123[0][0] ;
 wire \as2650.r123[0][1] ;
 wire \as2650.r123[0][2] ;
 wire \as2650.r123[0][3] ;
 wire \as2650.r123[0][4] ;
 wire \as2650.r123[0][5] ;
 wire \as2650.r123[0][6] ;
 wire \as2650.r123[0][7] ;
 wire \as2650.r123[1][0] ;
 wire \as2650.r123[1][1] ;
 wire \as2650.r123[1][2] ;
 wire \as2650.r123[1][3] ;
 wire \as2650.r123[1][4] ;
 wire \as2650.r123[1][5] ;
 wire \as2650.r123[1][6] ;
 wire \as2650.r123[1][7] ;
 wire \as2650.r123[2][0] ;
 wire \as2650.r123[2][1] ;
 wire \as2650.r123[2][2] ;
 wire \as2650.r123[2][3] ;
 wire \as2650.r123[2][4] ;
 wire \as2650.r123[2][5] ;
 wire \as2650.r123[2][6] ;
 wire \as2650.r123[2][7] ;
 wire \as2650.r123[3][0] ;
 wire \as2650.r123[3][1] ;
 wire \as2650.r123[3][2] ;
 wire \as2650.r123[3][3] ;
 wire \as2650.r123[3][4] ;
 wire \as2650.r123[3][5] ;
 wire \as2650.r123[3][6] ;
 wire \as2650.r123[3][7] ;
 wire \as2650.r123_2[0][0] ;
 wire \as2650.r123_2[0][1] ;
 wire \as2650.r123_2[0][2] ;
 wire \as2650.r123_2[0][3] ;
 wire \as2650.r123_2[0][4] ;
 wire \as2650.r123_2[0][5] ;
 wire \as2650.r123_2[0][6] ;
 wire \as2650.r123_2[0][7] ;
 wire \as2650.r123_2[1][0] ;
 wire \as2650.r123_2[1][1] ;
 wire \as2650.r123_2[1][2] ;
 wire \as2650.r123_2[1][3] ;
 wire \as2650.r123_2[1][4] ;
 wire \as2650.r123_2[1][5] ;
 wire \as2650.r123_2[1][6] ;
 wire \as2650.r123_2[1][7] ;
 wire \as2650.r123_2[2][0] ;
 wire \as2650.r123_2[2][1] ;
 wire \as2650.r123_2[2][2] ;
 wire \as2650.r123_2[2][3] ;
 wire \as2650.r123_2[2][4] ;
 wire \as2650.r123_2[2][5] ;
 wire \as2650.r123_2[2][6] ;
 wire \as2650.r123_2[2][7] ;
 wire \as2650.stack[0][0] ;
 wire \as2650.stack[0][10] ;
 wire \as2650.stack[0][11] ;
 wire \as2650.stack[0][12] ;
 wire \as2650.stack[0][1] ;
 wire \as2650.stack[0][2] ;
 wire \as2650.stack[0][3] ;
 wire \as2650.stack[0][4] ;
 wire \as2650.stack[0][5] ;
 wire \as2650.stack[0][6] ;
 wire \as2650.stack[0][7] ;
 wire \as2650.stack[0][8] ;
 wire \as2650.stack[0][9] ;
 wire \as2650.stack[1][0] ;
 wire \as2650.stack[1][10] ;
 wire \as2650.stack[1][11] ;
 wire \as2650.stack[1][12] ;
 wire \as2650.stack[1][1] ;
 wire \as2650.stack[1][2] ;
 wire \as2650.stack[1][3] ;
 wire \as2650.stack[1][4] ;
 wire \as2650.stack[1][5] ;
 wire \as2650.stack[1][6] ;
 wire \as2650.stack[1][7] ;
 wire \as2650.stack[1][8] ;
 wire \as2650.stack[1][9] ;
 wire \as2650.stack[2][0] ;
 wire \as2650.stack[2][10] ;
 wire \as2650.stack[2][11] ;
 wire \as2650.stack[2][12] ;
 wire \as2650.stack[2][1] ;
 wire \as2650.stack[2][2] ;
 wire \as2650.stack[2][3] ;
 wire \as2650.stack[2][4] ;
 wire \as2650.stack[2][5] ;
 wire \as2650.stack[2][6] ;
 wire \as2650.stack[2][7] ;
 wire \as2650.stack[2][8] ;
 wire \as2650.stack[2][9] ;
 wire \as2650.stack[3][0] ;
 wire \as2650.stack[3][10] ;
 wire \as2650.stack[3][11] ;
 wire \as2650.stack[3][12] ;
 wire \as2650.stack[3][1] ;
 wire \as2650.stack[3][2] ;
 wire \as2650.stack[3][3] ;
 wire \as2650.stack[3][4] ;
 wire \as2650.stack[3][5] ;
 wire \as2650.stack[3][6] ;
 wire \as2650.stack[3][7] ;
 wire \as2650.stack[3][8] ;
 wire \as2650.stack[3][9] ;
 wire \as2650.stack[4][0] ;
 wire \as2650.stack[4][10] ;
 wire \as2650.stack[4][11] ;
 wire \as2650.stack[4][12] ;
 wire \as2650.stack[4][1] ;
 wire \as2650.stack[4][2] ;
 wire \as2650.stack[4][3] ;
 wire \as2650.stack[4][4] ;
 wire \as2650.stack[4][5] ;
 wire \as2650.stack[4][6] ;
 wire \as2650.stack[4][7] ;
 wire \as2650.stack[4][8] ;
 wire \as2650.stack[4][9] ;
 wire \as2650.stack[5][0] ;
 wire \as2650.stack[5][10] ;
 wire \as2650.stack[5][11] ;
 wire \as2650.stack[5][12] ;
 wire \as2650.stack[5][1] ;
 wire \as2650.stack[5][2] ;
 wire \as2650.stack[5][3] ;
 wire \as2650.stack[5][4] ;
 wire \as2650.stack[5][5] ;
 wire \as2650.stack[5][6] ;
 wire \as2650.stack[5][7] ;
 wire \as2650.stack[5][8] ;
 wire \as2650.stack[5][9] ;
 wire \as2650.stack[6][0] ;
 wire \as2650.stack[6][10] ;
 wire \as2650.stack[6][11] ;
 wire \as2650.stack[6][12] ;
 wire \as2650.stack[6][1] ;
 wire \as2650.stack[6][2] ;
 wire \as2650.stack[6][3] ;
 wire \as2650.stack[6][4] ;
 wire \as2650.stack[6][5] ;
 wire \as2650.stack[6][6] ;
 wire \as2650.stack[6][7] ;
 wire \as2650.stack[6][8] ;
 wire \as2650.stack[6][9] ;
 wire \as2650.stack[7][0] ;
 wire \as2650.stack[7][10] ;
 wire \as2650.stack[7][11] ;
 wire \as2650.stack[7][12] ;
 wire \as2650.stack[7][1] ;
 wire \as2650.stack[7][2] ;
 wire \as2650.stack[7][3] ;
 wire \as2650.stack[7][4] ;
 wire \as2650.stack[7][5] ;
 wire \as2650.stack[7][6] ;
 wire \as2650.stack[7][7] ;
 wire \as2650.stack[7][8] ;
 wire \as2650.stack[7][9] ;
 wire \as2650.stack_ptr[0] ;
 wire \as2650.stack_ptr[1] ;
 wire \as2650.stack_ptr[2] ;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire clknet_leaf_0_wb_clk_i;
 wire net54;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net83;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire clknet_leaf_1_wb_clk_i;
 wire clknet_leaf_2_wb_clk_i;
 wire clknet_leaf_3_wb_clk_i;
 wire clknet_leaf_4_wb_clk_i;
 wire clknet_leaf_6_wb_clk_i;
 wire clknet_leaf_7_wb_clk_i;
 wire clknet_leaf_8_wb_clk_i;
 wire clknet_leaf_9_wb_clk_i;
 wire clknet_leaf_10_wb_clk_i;
 wire clknet_leaf_12_wb_clk_i;
 wire clknet_leaf_13_wb_clk_i;
 wire clknet_leaf_14_wb_clk_i;
 wire clknet_leaf_15_wb_clk_i;
 wire clknet_leaf_16_wb_clk_i;
 wire clknet_leaf_17_wb_clk_i;
 wire clknet_leaf_19_wb_clk_i;
 wire clknet_leaf_21_wb_clk_i;
 wire clknet_leaf_24_wb_clk_i;
 wire clknet_leaf_25_wb_clk_i;
 wire clknet_leaf_27_wb_clk_i;
 wire clknet_leaf_28_wb_clk_i;
 wire clknet_leaf_29_wb_clk_i;
 wire clknet_leaf_30_wb_clk_i;
 wire clknet_leaf_31_wb_clk_i;
 wire clknet_leaf_32_wb_clk_i;
 wire clknet_leaf_33_wb_clk_i;
 wire clknet_leaf_34_wb_clk_i;
 wire clknet_leaf_35_wb_clk_i;
 wire clknet_leaf_36_wb_clk_i;
 wire clknet_leaf_37_wb_clk_i;
 wire clknet_leaf_38_wb_clk_i;
 wire clknet_leaf_39_wb_clk_i;
 wire clknet_leaf_40_wb_clk_i;
 wire clknet_leaf_41_wb_clk_i;
 wire clknet_leaf_42_wb_clk_i;
 wire clknet_leaf_43_wb_clk_i;
 wire clknet_leaf_44_wb_clk_i;
 wire clknet_leaf_45_wb_clk_i;
 wire clknet_leaf_46_wb_clk_i;
 wire clknet_leaf_47_wb_clk_i;
 wire clknet_leaf_48_wb_clk_i;
 wire clknet_leaf_49_wb_clk_i;
 wire clknet_leaf_50_wb_clk_i;
 wire clknet_leaf_51_wb_clk_i;
 wire clknet_leaf_52_wb_clk_i;
 wire clknet_leaf_53_wb_clk_i;
 wire clknet_leaf_54_wb_clk_i;
 wire clknet_leaf_55_wb_clk_i;
 wire clknet_leaf_56_wb_clk_i;
 wire clknet_leaf_57_wb_clk_i;
 wire clknet_leaf_60_wb_clk_i;
 wire clknet_leaf_61_wb_clk_i;
 wire clknet_leaf_62_wb_clk_i;
 wire clknet_leaf_63_wb_clk_i;
 wire clknet_leaf_64_wb_clk_i;
 wire clknet_leaf_65_wb_clk_i;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0_0_wb_clk_i;
 wire clknet_3_1_0_wb_clk_i;
 wire clknet_3_2_0_wb_clk_i;
 wire clknet_3_3_0_wb_clk_i;
 wire clknet_3_4_0_wb_clk_i;
 wire clknet_3_5_0_wb_clk_i;
 wire clknet_3_6_0_wb_clk_i;
 wire clknet_3_7_0_wb_clk_i;
 wire clknet_opt_1_0_wb_clk_i;
 wire clknet_opt_2_0_wb_clk_i;
 wire clknet_opt_2_1_wb_clk_i;
 wire clknet_opt_3_0_wb_clk_i;
 wire clknet_opt_3_1_wb_clk_i;
 wire clknet_opt_4_0_wb_clk_i;

 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3594_ (.I(net23),
    .ZN(net18));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3595_ (.I(\as2650.ins_reg[1] ),
    .Z(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3596_ (.I(_3131_),
    .ZN(_3132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3597_ (.I(_3132_),
    .Z(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3598_ (.I(\as2650.ins_reg[0] ),
    .ZN(_3134_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3599_ (.I(_3134_),
    .Z(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3600_ (.A1(_3133_),
    .A2(_3135_),
    .ZN(_3136_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3601_ (.I(_3136_),
    .Z(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3602_ (.I(_3137_),
    .Z(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3603_ (.A1(\as2650.halted ),
    .A2(net10),
    .ZN(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3604_ (.I(_3139_),
    .Z(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3605_ (.I(\as2650.cycle[7] ),
    .ZN(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3606_ (.A1(\as2650.cycle[5] ),
    .A2(\as2650.cycle[4] ),
    .ZN(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3607_ (.A1(_3141_),
    .A2(_3142_),
    .ZN(_3143_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3608_ (.A1(\as2650.cycle[6] ),
    .A2(_3143_),
    .ZN(_3144_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3609_ (.A1(\as2650.cycle[3] ),
    .A2(\as2650.cycle[2] ),
    .ZN(_3145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3610_ (.A1(_3144_),
    .A2(_3145_),
    .ZN(_3146_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3611_ (.I(_3146_),
    .Z(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3612_ (.I(\as2650.cycle[0] ),
    .ZN(_3148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3613_ (.A1(\as2650.cycle[1] ),
    .A2(_3148_),
    .ZN(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3614_ (.A1(_3147_),
    .A2(_3149_),
    .ZN(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3615_ (.I(_3150_),
    .Z(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3616_ (.I(_3151_),
    .Z(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3617_ (.I(\as2650.ins_reg[3] ),
    .Z(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3618_ (.I(_3153_),
    .Z(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3619_ (.I(\as2650.ins_reg[2] ),
    .Z(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3620_ (.I(_3155_),
    .Z(_3156_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3621_ (.I(_3156_),
    .ZN(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3622_ (.I(\as2650.ins_reg[4] ),
    .Z(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3623_ (.I(\as2650.ins_reg[5] ),
    .Z(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3624_ (.I(_3159_),
    .Z(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3625_ (.I(\as2650.ins_reg[6] ),
    .Z(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3626_ (.I(\as2650.ins_reg[7] ),
    .Z(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3627_ (.I(_3162_),
    .ZN(_3163_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3628_ (.A1(_3161_),
    .A2(_3163_),
    .ZN(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3629_ (.A1(_3160_),
    .A2(_3164_),
    .ZN(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3630_ (.A1(_3157_),
    .A2(_3158_),
    .A3(_3165_),
    .ZN(_3166_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3631_ (.A1(_3154_),
    .A2(_3166_),
    .ZN(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3632_ (.I(_3167_),
    .Z(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3633_ (.I(_3154_),
    .Z(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3634_ (.I(\as2650.ins_reg[4] ),
    .Z(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3635_ (.I(_3170_),
    .Z(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3636_ (.I(_3171_),
    .Z(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3637_ (.I(_3161_),
    .Z(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3638_ (.I(_3173_),
    .Z(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3639_ (.I(_3150_),
    .Z(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3640_ (.I(_3175_),
    .Z(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3641_ (.A1(_3169_),
    .A2(_3172_),
    .A3(_3174_),
    .A4(_3176_),
    .ZN(_3177_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3642_ (.I(_3170_),
    .ZN(_3178_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3643_ (.I(_3178_),
    .Z(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3644_ (.I(\as2650.cycle[1] ),
    .ZN(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3645_ (.I(\as2650.cycle[0] ),
    .Z(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3646_ (.A1(_3180_),
    .A2(_3181_),
    .ZN(_3182_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3647_ (.A1(\as2650.cycle[6] ),
    .A2(_3145_),
    .ZN(_3183_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _3648_ (.A1(_3143_),
    .A2(_3182_),
    .A3(_3183_),
    .ZN(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3649_ (.I(\as2650.idx_ctrl[1] ),
    .ZN(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3650_ (.I(\as2650.idx_ctrl[0] ),
    .ZN(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3651_ (.A1(_3185_),
    .A2(_3186_),
    .ZN(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3652_ (.A1(_3179_),
    .A2(_3184_),
    .A3(_3187_),
    .ZN(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3653_ (.A1(_3177_),
    .A2(_3188_),
    .ZN(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3654_ (.A1(_3152_),
    .A2(_3168_),
    .B(_3189_),
    .ZN(_3190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3655_ (.I(\as2650.psl[4] ),
    .Z(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3656_ (.I(_3191_),
    .Z(_3192_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3657_ (.I(_3192_),
    .Z(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3658_ (.I(_3193_),
    .Z(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3659_ (.I(_3194_),
    .Z(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3660_ (.I(\as2650.ins_reg[1] ),
    .Z(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3661_ (.I(_3196_),
    .Z(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3662_ (.I(\as2650.ins_reg[0] ),
    .Z(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3663_ (.A1(_3197_),
    .A2(_3198_),
    .ZN(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3664_ (.I(_3199_),
    .Z(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3665_ (.A1(_3195_),
    .A2(_3200_),
    .Z(_3201_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3666_ (.I(_3153_),
    .ZN(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3667_ (.I(_3202_),
    .Z(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3668_ (.I(_3203_),
    .Z(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3669_ (.A1(_3195_),
    .A2(_3200_),
    .ZN(_3205_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3670_ (.I(_3155_),
    .Z(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3671_ (.I(_3206_),
    .Z(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3672_ (.I(_3162_),
    .Z(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3673_ (.I(_3208_),
    .Z(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3674_ (.A1(_3158_),
    .A2(_3160_),
    .ZN(_3210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3675_ (.I(_3210_),
    .Z(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3676_ (.A1(_3207_),
    .A2(_3209_),
    .A3(_3211_),
    .ZN(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3677_ (.I(_3144_),
    .Z(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3678_ (.I(_3213_),
    .Z(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3679_ (.I(\as2650.cycle[3] ),
    .Z(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3680_ (.I(\as2650.cycle[2] ),
    .Z(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3681_ (.I(_3216_),
    .Z(_3217_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3682_ (.I(\as2650.cycle[1] ),
    .Z(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3683_ (.A1(_3218_),
    .A2(\as2650.cycle[0] ),
    .ZN(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _3684_ (.A1(_3215_),
    .A2(_3217_),
    .A3(_3219_),
    .ZN(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3685_ (.A1(_3214_),
    .A2(_3220_),
    .Z(_3221_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3686_ (.I(_3221_),
    .Z(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _3687_ (.A1(_3204_),
    .A2(_3205_),
    .A3(_3212_),
    .A4(_3222_),
    .ZN(_3223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3688_ (.I(\as2650.cycle[7] ),
    .Z(_3224_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3689_ (.A1(_3224_),
    .A2(_3142_),
    .ZN(_3225_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3690_ (.A1(_3182_),
    .A2(_3183_),
    .A3(_3225_),
    .Z(_3226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3691_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3226_),
    .ZN(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3692_ (.I(\as2650.addr_buff[5] ),
    .Z(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3693_ (.I(\as2650.addr_buff[6] ),
    .Z(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3694_ (.A1(_3228_),
    .A2(_3229_),
    .ZN(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3695_ (.A1(_3172_),
    .A2(_3230_),
    .ZN(_3231_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3696_ (.I(_3231_),
    .Z(_3232_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3697_ (.A1(_3205_),
    .A2(_3227_),
    .A3(_3232_),
    .ZN(_3233_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3698_ (.A1(_3190_),
    .A2(_3201_),
    .B(_3223_),
    .C(_3233_),
    .ZN(_3234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3699_ (.A1(_3140_),
    .A2(_3234_),
    .ZN(_3235_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3700_ (.I(_3152_),
    .Z(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3701_ (.I(\as2650.halted ),
    .ZN(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3702_ (.I(net10),
    .ZN(_3238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3703_ (.A1(_3237_),
    .A2(_3238_),
    .ZN(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3704_ (.A1(_3239_),
    .A2(_3201_),
    .ZN(_3240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3705_ (.I(_3240_),
    .Z(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3706_ (.A1(\as2650.ins_reg[6] ),
    .A2(\as2650.ins_reg[7] ),
    .ZN(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3707_ (.A1(_3159_),
    .A2(_3242_),
    .ZN(_3243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3708_ (.I(_3243_),
    .Z(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3709_ (.A1(\as2650.ins_reg[2] ),
    .A2(\as2650.ins_reg[3] ),
    .Z(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3710_ (.I(_3245_),
    .Z(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3711_ (.I(_3246_),
    .Z(_3247_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3712_ (.I(_3247_),
    .Z(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3713_ (.A1(_3171_),
    .A2(_3248_),
    .ZN(_3249_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3714_ (.I(_3249_),
    .Z(_3250_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3715_ (.A1(_3244_),
    .A2(_3250_),
    .Z(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3716_ (.A1(_3236_),
    .A2(_3241_),
    .A3(_3251_),
    .ZN(_3252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3717_ (.I(_3195_),
    .Z(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3718_ (.I(_3158_),
    .Z(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3719_ (.I(_3254_),
    .Z(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3720_ (.I(_3255_),
    .Z(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3721_ (.A1(_3155_),
    .A2(_3153_),
    .ZN(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3722_ (.I(_3257_),
    .Z(_3258_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3723_ (.I(_3258_),
    .Z(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3724_ (.I(_3259_),
    .Z(_3260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3725_ (.I(_3260_),
    .Z(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3726_ (.I(_3200_),
    .Z(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3727_ (.I(\as2650.ins_reg[5] ),
    .ZN(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3728_ (.A1(_3263_),
    .A2(_3242_),
    .ZN(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _3729_ (.A1(_3261_),
    .A2(_3187_),
    .A3(_3262_),
    .A4(_3264_),
    .ZN(_3265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3730_ (.I(_3218_),
    .Z(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3731_ (.I(\as2650.cycle[3] ),
    .ZN(_3267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3732_ (.I(_3267_),
    .Z(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3733_ (.A1(_3268_),
    .A2(_3217_),
    .A3(_3213_),
    .ZN(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3734_ (.A1(_3266_),
    .A2(_3181_),
    .A3(_3269_),
    .ZN(_3270_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3735_ (.I(_3270_),
    .Z(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3736_ (.A1(_3265_),
    .A2(_3271_),
    .ZN(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _3737_ (.A1(_3253_),
    .A2(_3256_),
    .A3(_3239_),
    .A4(_3272_),
    .Z(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3738_ (.I(_3148_),
    .Z(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3739_ (.A1(_3180_),
    .A2(_3146_),
    .ZN(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3740_ (.A1(_3274_),
    .A2(_3275_),
    .ZN(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3741_ (.A1(_3139_),
    .A2(_3205_),
    .ZN(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3742_ (.A1(_3276_),
    .A2(_3277_),
    .ZN(_3278_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3743_ (.I(_3153_),
    .Z(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3744_ (.A1(\as2650.ins_reg[4] ),
    .A2(\as2650.ins_reg[6] ),
    .A3(_3162_),
    .ZN(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3745_ (.A1(_3159_),
    .A2(_3280_),
    .ZN(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3746_ (.I(_3281_),
    .Z(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3747_ (.A1(_3157_),
    .A2(_3282_),
    .ZN(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3748_ (.A1(_3279_),
    .A2(_3283_),
    .ZN(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3749_ (.I(_3284_),
    .Z(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3750_ (.A1(_3278_),
    .A2(_3285_),
    .ZN(_3286_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _3751_ (.A1(_3235_),
    .A2(_3252_),
    .A3(_3273_),
    .A4(_3286_),
    .ZN(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3752_ (.I(_3287_),
    .Z(_3288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3753_ (.A1(_3138_),
    .A2(_3288_),
    .ZN(_3289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3754_ (.I(_3289_),
    .Z(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3755_ (.I0(\as2650.r123[0][0] ),
    .I1(\as2650.r123_2[0][0] ),
    .S(\as2650.psl[4] ),
    .Z(_3291_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3756_ (.I0(\as2650.r123[1][0] ),
    .I1(\as2650.r123_2[1][0] ),
    .S(\as2650.psl[4] ),
    .Z(_3292_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3757_ (.I0(\as2650.r123[2][0] ),
    .I1(\as2650.r123_2[2][0] ),
    .S(\as2650.psl[4] ),
    .Z(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3758_ (.I0(\as2650.r0[0] ),
    .I1(_3291_),
    .I2(_3292_),
    .I3(_3293_),
    .S0(\as2650.ins_reg[0] ),
    .S1(_3131_),
    .Z(_3294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3759_ (.I(_3294_),
    .Z(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _3760_ (.I(_3295_),
    .ZN(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3761_ (.I(_3296_),
    .Z(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3762_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3186_),
    .ZN(_3298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3763_ (.A1(_3185_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_3299_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3764_ (.A1(_3298_),
    .A2(_3299_),
    .ZN(_3300_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3765_ (.A1(_3297_),
    .A2(_3300_),
    .Z(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3766_ (.I(_3301_),
    .Z(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3767_ (.I(_3255_),
    .Z(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3768_ (.I(_3182_),
    .Z(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _3769_ (.A1(_3143_),
    .A2(_3304_),
    .A3(_3183_),
    .Z(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3770_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_3306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3771_ (.I(_3306_),
    .Z(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3772_ (.A1(_3303_),
    .A2(_3305_),
    .A3(_3307_),
    .ZN(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3773_ (.A1(_3308_),
    .A2(_3241_),
    .ZN(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3774_ (.I(_3309_),
    .Z(_3310_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3775_ (.I(\as2650.r0[0] ),
    .Z(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3776_ (.A1(_3251_),
    .A2(_3278_),
    .ZN(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3777_ (.I(_3312_),
    .Z(_3313_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3778_ (.I(_3227_),
    .Z(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _3779_ (.A1(_3241_),
    .A2(_3314_),
    .A3(_3232_),
    .ZN(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3780_ (.I(_3175_),
    .Z(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3781_ (.A1(_3316_),
    .A2(_3241_),
    .A3(_3284_),
    .ZN(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3782_ (.I(_3317_),
    .Z(_3318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3783_ (.I(\as2650.psl[3] ),
    .Z(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3784_ (.A1(\as2650.r0[7] ),
    .A2(_3199_),
    .ZN(_3320_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3785_ (.I0(\as2650.r123[2][7] ),
    .I1(\as2650.r123_2[2][7] ),
    .S(_3193_),
    .Z(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3786_ (.A1(_3137_),
    .A2(_3321_),
    .ZN(_3322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3787_ (.I(_3191_),
    .Z(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3788_ (.I(_3323_),
    .Z(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3789_ (.I(_3324_),
    .Z(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3790_ (.A1(_3133_),
    .A2(_3198_),
    .ZN(_3326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3791_ (.I(_3326_),
    .Z(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3792_ (.I(\as2650.r123_2[1][7] ),
    .ZN(_3328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3793_ (.A1(_3325_),
    .A2(_3328_),
    .ZN(_3329_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3794_ (.A1(_3325_),
    .A2(\as2650.r123[1][7] ),
    .B(_3327_),
    .C(_3329_),
    .ZN(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3795_ (.I(_3131_),
    .Z(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3796_ (.I(_3134_),
    .Z(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3797_ (.A1(_3331_),
    .A2(_3332_),
    .ZN(_3333_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3798_ (.I(\as2650.r123_2[0][7] ),
    .ZN(_3334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3799_ (.A1(_3325_),
    .A2(_3334_),
    .ZN(_3335_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _3800_ (.A1(_3194_),
    .A2(\as2650.r123[0][7] ),
    .B(_3333_),
    .C(_3335_),
    .ZN(_3336_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _3801_ (.A1(_3320_),
    .A2(_3322_),
    .A3(_3330_),
    .A4(_3336_),
    .Z(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3802_ (.I(_3337_),
    .Z(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3803_ (.I(_3338_),
    .Z(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3804_ (.I(_3339_),
    .Z(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3805_ (.A1(\as2650.psl[3] ),
    .A2(\as2650.carry ),
    .ZN(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3806_ (.A1(_3319_),
    .A2(_3340_),
    .B(_3341_),
    .ZN(_3342_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3807_ (.I(_3342_),
    .ZN(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3808_ (.A1(_3168_),
    .A2(_3278_),
    .ZN(_3344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3809_ (.I(_3344_),
    .Z(_3345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3810_ (.I(\as2650.ins_reg[0] ),
    .Z(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3811_ (.I0(\as2650.r123[0][1] ),
    .I1(\as2650.r123[2][1] ),
    .I2(\as2650.r123_2[0][1] ),
    .I3(\as2650.r123_2[2][1] ),
    .S0(_3196_),
    .S1(_3323_),
    .Z(_3347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3812_ (.A1(_3346_),
    .A2(_3347_),
    .ZN(_3348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3813_ (.I(_3191_),
    .Z(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3814_ (.I0(\as2650.r123[1][1] ),
    .I1(\as2650.r123_2[1][1] ),
    .S(_3349_),
    .Z(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3815_ (.A1(\as2650.r0[1] ),
    .A2(_3331_),
    .Z(_3351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3816_ (.A1(_3133_),
    .A2(_3350_),
    .B(_3351_),
    .C(_3332_),
    .ZN(_3352_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3817_ (.A1(_3348_),
    .A2(_3352_),
    .ZN(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3818_ (.I(_3353_),
    .Z(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3819_ (.I(_3354_),
    .Z(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3820_ (.I(_3163_),
    .Z(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3821_ (.A1(_3156_),
    .A2(_3210_),
    .ZN(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3822_ (.A1(_3356_),
    .A2(_3357_),
    .ZN(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3823_ (.A1(_3144_),
    .A2(_3145_),
    .Z(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3824_ (.A1(_3180_),
    .A2(_3148_),
    .ZN(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3825_ (.A1(_3359_),
    .A2(_3360_),
    .ZN(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3826_ (.I(_3361_),
    .Z(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _3827_ (.A1(_3154_),
    .A2(_3358_),
    .A3(_3362_),
    .ZN(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3828_ (.A1(_3240_),
    .A2(_3363_),
    .ZN(_3364_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3829_ (.I(_3364_),
    .ZN(_3365_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3830_ (.I(_3365_),
    .Z(_3366_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3831_ (.I(_3295_),
    .Z(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3832_ (.I(_3367_),
    .Z(_3368_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3833_ (.I(_3368_),
    .Z(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3834_ (.A1(_3280_),
    .A2(_3369_),
    .Z(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3835_ (.I(_3344_),
    .Z(_3371_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3836_ (.I(net1),
    .Z(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3837_ (.I(_3372_),
    .Z(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3838_ (.I(_3373_),
    .Z(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3839_ (.A1(_3374_),
    .A2(_3365_),
    .ZN(_3375_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3840_ (.A1(_3366_),
    .A2(_3370_),
    .B(_3371_),
    .C(_3375_),
    .ZN(_3376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3841_ (.I(_3317_),
    .Z(_3377_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3842_ (.A1(_3345_),
    .A2(_3355_),
    .B(_3376_),
    .C(_3377_),
    .ZN(_3378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3843_ (.I(_3312_),
    .Z(_3379_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3844_ (.A1(_3318_),
    .A2(_3343_),
    .B(_3378_),
    .C(_3379_),
    .ZN(_3380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3845_ (.A1(_3311_),
    .A2(_3313_),
    .B(_3315_),
    .C(_3380_),
    .ZN(_3381_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3846_ (.A1(_3227_),
    .A2(_3231_),
    .ZN(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3847_ (.A1(_3277_),
    .A2(_3382_),
    .ZN(_3383_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3848_ (.I(_3383_),
    .Z(_3384_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3849_ (.I(\as2650.addr_buff[5] ),
    .ZN(_3385_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3850_ (.A1(_3385_),
    .A2(\as2650.addr_buff[6] ),
    .ZN(_3386_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3851_ (.I(\as2650.addr_buff[6] ),
    .ZN(_3387_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3852_ (.A1(\as2650.addr_buff[5] ),
    .A2(_3387_),
    .ZN(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_4 _3853_ (.A1(_3386_),
    .A2(_3388_),
    .ZN(_3389_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3854_ (.A1(_3297_),
    .A2(_3389_),
    .Z(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3855_ (.I(_3390_),
    .Z(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3856_ (.A1(_3384_),
    .A2(_3391_),
    .ZN(_3392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3857_ (.A1(_3381_),
    .A2(_3392_),
    .A3(_3310_),
    .ZN(_3393_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3858_ (.A1(_3302_),
    .A2(_3310_),
    .B(_3393_),
    .ZN(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3859_ (.I(_3160_),
    .Z(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3860_ (.A1(_3161_),
    .A2(_3208_),
    .ZN(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3861_ (.A1(_3395_),
    .A2(_3396_),
    .Z(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3862_ (.I(_3397_),
    .Z(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3863_ (.I0(\as2650.holding_reg[0] ),
    .I1(_3294_),
    .S(_3246_),
    .Z(_3399_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3864_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3245_),
    .Z(_3400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _3865_ (.A1(_3257_),
    .A2(_3295_),
    .B(_3400_),
    .ZN(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3866_ (.A1(_3399_),
    .A2(_3401_),
    .ZN(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3867_ (.I(_3341_),
    .ZN(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3868_ (.I(_3263_),
    .Z(_3404_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3869_ (.A1(_3161_),
    .A2(_3163_),
    .ZN(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3870_ (.I(_3405_),
    .Z(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3871_ (.A1(_3404_),
    .A2(_3406_),
    .ZN(_3407_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3872_ (.I(_3407_),
    .Z(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3873_ (.A1(_3403_),
    .A2(_3402_),
    .B(_3408_),
    .ZN(_3409_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3874_ (.A1(_3403_),
    .A2(_3402_),
    .B(_3409_),
    .ZN(_3410_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3875_ (.I(\as2650.carry ),
    .ZN(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3876_ (.A1(\as2650.psl[3] ),
    .A2(_3411_),
    .ZN(_3412_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3877_ (.A1(_3399_),
    .A2(_3401_),
    .Z(_3413_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3878_ (.I(_3413_),
    .Z(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3879_ (.A1(_3395_),
    .A2(_3406_),
    .ZN(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3880_ (.A1(_3412_),
    .A2(_3414_),
    .B(_3415_),
    .ZN(_3416_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3881_ (.A1(_3412_),
    .A2(_3414_),
    .B(_3416_),
    .ZN(_3417_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _3882_ (.I(\as2650.ins_reg[6] ),
    .ZN(_3418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3883_ (.A1(_3418_),
    .A2(_3162_),
    .ZN(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3884_ (.I(_3419_),
    .Z(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3885_ (.I(_3399_),
    .Z(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3886_ (.A1(_3263_),
    .A2(_3419_),
    .ZN(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3887_ (.I(_3422_),
    .Z(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3888_ (.A1(_3401_),
    .A2(_3406_),
    .B(_3423_),
    .ZN(_3424_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3889_ (.A1(_3420_),
    .A2(_3421_),
    .B(_3424_),
    .ZN(_3425_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _3890_ (.A1(_3410_),
    .A2(_3417_),
    .A3(_3425_),
    .ZN(_3426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3891_ (.A1(\as2650.holding_reg[0] ),
    .A2(_3367_),
    .ZN(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3892_ (.I(_3397_),
    .Z(_3428_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3893_ (.A1(_3165_),
    .A2(_3427_),
    .B(_3428_),
    .ZN(_3429_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _3894_ (.A1(_3398_),
    .A2(_3402_),
    .B1(_3426_),
    .B2(_3429_),
    .ZN(_3430_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3895_ (.I(_3430_),
    .Z(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3896_ (.I(_3253_),
    .Z(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3897_ (.I(_3303_),
    .Z(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3898_ (.I(_3239_),
    .Z(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _3899_ (.A1(_3432_),
    .A2(_3433_),
    .A3(_3434_),
    .A4(_3272_),
    .ZN(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3900_ (.I(_3435_),
    .Z(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3901_ (.I0(_3394_),
    .I1(_3431_),
    .S(_3436_),
    .Z(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3902_ (.I(net10),
    .Z(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3903_ (.A1(_3138_),
    .A2(_3287_),
    .B(_3438_),
    .ZN(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3904_ (.I(_3439_),
    .Z(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3905_ (.A1(\as2650.r123[2][0] ),
    .A2(_3440_),
    .ZN(_3441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3906_ (.A1(_3290_),
    .A2(_3437_),
    .B(_3441_),
    .ZN(_0000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3907_ (.A1(_3188_),
    .A2(_3277_),
    .ZN(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3908_ (.I(_3442_),
    .Z(_3443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3909_ (.I(_3383_),
    .Z(_3444_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3910_ (.I(_3353_),
    .Z(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3911_ (.A1(\as2650.addr_buff[5] ),
    .A2(_3387_),
    .ZN(_3446_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3912_ (.A1(_3367_),
    .A2(_3446_),
    .B(_3388_),
    .ZN(_3447_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3913_ (.A1(_3296_),
    .A2(_3445_),
    .A3(_3447_),
    .Z(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3914_ (.I(_3448_),
    .Z(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3915_ (.I(_3317_),
    .Z(_3450_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3916_ (.I(_3369_),
    .Z(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3917_ (.I(_3344_),
    .Z(_3452_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3918_ (.I0(\as2650.r123[1][2] ),
    .I1(\as2650.r123_2[1][2] ),
    .S(_3191_),
    .Z(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3919_ (.A1(\as2650.r0[2] ),
    .A2(_3196_),
    .Z(_3454_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3920_ (.A1(_3132_),
    .A2(_3453_),
    .B(_3454_),
    .C(_3332_),
    .ZN(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3921_ (.I0(\as2650.r123[0][2] ),
    .I1(\as2650.r123[2][2] ),
    .I2(\as2650.r123_2[0][2] ),
    .I3(\as2650.r123_2[2][2] ),
    .S0(_3131_),
    .S1(_3349_),
    .Z(_3456_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3922_ (.A1(_3198_),
    .A2(_3456_),
    .ZN(_3457_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3923_ (.A1(_3455_),
    .A2(_3457_),
    .Z(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3924_ (.I(_3458_),
    .Z(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3925_ (.I(_3459_),
    .Z(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3926_ (.I(_3460_),
    .Z(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3927_ (.I(net2),
    .Z(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3928_ (.I(_3462_),
    .Z(_3463_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3929_ (.I(_3463_),
    .Z(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3930_ (.I(_3464_),
    .Z(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3931_ (.I(_3465_),
    .Z(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3932_ (.I(_3364_),
    .Z(_3467_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3933_ (.I(_3344_),
    .Z(_3468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3934_ (.I(_3364_),
    .Z(_3469_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3935_ (.A1(_3348_),
    .A2(_3352_),
    .Z(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3936_ (.I(_3470_),
    .Z(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3937_ (.I(_3471_),
    .Z(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3938_ (.A1(\as2650.ins_reg[4] ),
    .A2(_3264_),
    .ZN(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3939_ (.A1(_3281_),
    .A2(_3368_),
    .ZN(_3474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3940_ (.A1(_3369_),
    .A2(_3473_),
    .B(_3474_),
    .ZN(_3475_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3941_ (.A1(_3472_),
    .A2(_3475_),
    .Z(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3942_ (.A1(_3469_),
    .A2(_3476_),
    .ZN(_3477_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3943_ (.A1(_3466_),
    .A2(_3467_),
    .B(_3468_),
    .C(_3477_),
    .ZN(_3478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3944_ (.I(_3317_),
    .Z(_3479_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3945_ (.A1(_3452_),
    .A2(_3461_),
    .B(_3478_),
    .C(_3479_),
    .ZN(_3480_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3946_ (.A1(_3450_),
    .A2(_3451_),
    .B(_3480_),
    .ZN(_3481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3947_ (.I(\as2650.r0[1] ),
    .Z(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3948_ (.I(_3482_),
    .Z(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3949_ (.I(_3312_),
    .Z(_3484_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3950_ (.A1(_3483_),
    .A2(_3484_),
    .B(_3315_),
    .ZN(_3485_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3951_ (.A1(_3313_),
    .A2(_3481_),
    .B(_3485_),
    .ZN(_3486_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3952_ (.A1(_3444_),
    .A2(_3449_),
    .B(_3486_),
    .ZN(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3953_ (.I(_3442_),
    .Z(_3488_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3954_ (.A1(_3185_),
    .A2(\as2650.idx_ctrl[0] ),
    .ZN(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3955_ (.A1(_3367_),
    .A2(_3489_),
    .B(_3299_),
    .ZN(_3490_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _3956_ (.A1(_3296_),
    .A2(_3445_),
    .A3(_3490_),
    .Z(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3957_ (.I(_3491_),
    .Z(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3958_ (.A1(_3488_),
    .A2(_3492_),
    .ZN(_3493_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3959_ (.I(_3273_),
    .Z(_3494_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3960_ (.A1(_3443_),
    .A2(_3487_),
    .B(_3493_),
    .C(_3494_),
    .ZN(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3961_ (.I(_3435_),
    .Z(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3962_ (.I(\as2650.holding_reg[1] ),
    .Z(_3497_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3963_ (.A1(_3497_),
    .A2(_3257_),
    .ZN(_3498_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3964_ (.A1(_3258_),
    .A2(_3471_),
    .B(_3498_),
    .ZN(_3499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3965_ (.I(_3499_),
    .Z(_3500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3966_ (.A1(_3397_),
    .A2(_3500_),
    .ZN(_3501_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3967_ (.I(\as2650.holding_reg[1] ),
    .Z(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3968_ (.A1(_3502_),
    .A2(_3354_),
    .Z(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _3969_ (.I(_3418_),
    .Z(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _3970_ (.A1(_3504_),
    .A2(_3208_),
    .ZN(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _3971_ (.A1(_3404_),
    .A2(_3505_),
    .ZN(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3972_ (.A1(_3497_),
    .A2(_3471_),
    .Z(_3507_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3973_ (.I(_3507_),
    .Z(_3508_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _3974_ (.A1(_3399_),
    .A2(_3427_),
    .B1(_3413_),
    .B2(_3412_),
    .ZN(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3975_ (.A1(_3508_),
    .A2(_3509_),
    .Z(_3510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3976_ (.A1(_3506_),
    .A2(_3510_),
    .ZN(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3977_ (.A1(_3160_),
    .A2(_3505_),
    .ZN(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _3978_ (.A1(_3341_),
    .A2(_3414_),
    .B(_3427_),
    .ZN(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _3979_ (.A1(_3507_),
    .A2(_3513_),
    .Z(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3980_ (.A1(_3260_),
    .A2(_3355_),
    .ZN(_3515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _3981_ (.A1(_3502_),
    .A2(_3248_),
    .B(_3405_),
    .ZN(_3516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _3982_ (.A1(_3404_),
    .A2(_3164_),
    .ZN(_3517_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _3983_ (.A1(_3512_),
    .A2(_3514_),
    .B1(_3515_),
    .B2(_3516_),
    .C(_3517_),
    .ZN(_3518_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _3984_ (.A1(_3511_),
    .A2(_3518_),
    .Z(_3519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3985_ (.A1(_3502_),
    .A2(_3355_),
    .B(_3419_),
    .ZN(_3520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3986_ (.A1(_3422_),
    .A2(_3520_),
    .ZN(_3521_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _3987_ (.A1(_3422_),
    .A2(_3503_),
    .B1(_3519_),
    .B2(_3521_),
    .ZN(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _3988_ (.A1(_3501_),
    .A2(_3522_),
    .ZN(_3523_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _3989_ (.I(_3523_),
    .Z(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3990_ (.A1(_3496_),
    .A2(_3524_),
    .ZN(_3525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3991_ (.A1(_3495_),
    .A2(_3525_),
    .ZN(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _3992_ (.A1(\as2650.r123[2][1] ),
    .A2(_3440_),
    .ZN(_3527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _3993_ (.A1(_3290_),
    .A2(_3526_),
    .B(_3527_),
    .ZN(_0001_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3994_ (.I(\as2650.r0[2] ),
    .Z(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _3995_ (.I(_3472_),
    .Z(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _3996_ (.I0(\as2650.r123[1][3] ),
    .I1(\as2650.r123_2[1][3] ),
    .S(_3349_),
    .Z(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _3997_ (.A1(\as2650.r0[3] ),
    .A2(_3331_),
    .Z(_3531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _3998_ (.A1(_3132_),
    .A2(_3530_),
    .B(_3531_),
    .C(_3332_),
    .ZN(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _3999_ (.I0(\as2650.r123[0][3] ),
    .I1(\as2650.r123[2][3] ),
    .I2(\as2650.r123_2[0][3] ),
    .I3(\as2650.r123_2[2][3] ),
    .S0(_3196_),
    .S1(_3349_),
    .Z(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4000_ (.A1(_3198_),
    .A2(_3533_),
    .ZN(_3534_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4001_ (.A1(_3532_),
    .A2(_3534_),
    .ZN(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4002_ (.I(_3535_),
    .Z(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4003_ (.I(_3536_),
    .Z(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4004_ (.I(net3),
    .Z(_3538_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4005_ (.I(_3538_),
    .ZN(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4006_ (.I(_3539_),
    .Z(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4007_ (.I(_3540_),
    .Z(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4008_ (.I(_3541_),
    .Z(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4009_ (.I(_3542_),
    .Z(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4010_ (.A1(_3455_),
    .A2(_3457_),
    .ZN(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4011_ (.I(_3544_),
    .Z(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4012_ (.I(_3545_),
    .Z(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4013_ (.A1(_3170_),
    .A2(_3243_),
    .ZN(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4014_ (.I(_3297_),
    .Z(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4015_ (.A1(_3263_),
    .A2(_3280_),
    .ZN(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4016_ (.I0(_3482_),
    .I1(_3350_),
    .S(_3197_),
    .Z(_3550_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4017_ (.A1(_3346_),
    .A2(_3347_),
    .Z(_3551_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4018_ (.A1(_3135_),
    .A2(_3550_),
    .B(_3551_),
    .C(_3295_),
    .ZN(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4019_ (.I(_3552_),
    .Z(_3553_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4020_ (.A1(_3549_),
    .A2(_3553_),
    .ZN(_3554_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4021_ (.A1(_3547_),
    .A2(_3548_),
    .A3(_3472_),
    .B(_3554_),
    .ZN(_3555_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4022_ (.A1(_3546_),
    .A2(_3555_),
    .Z(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4023_ (.A1(_3469_),
    .A2(_3556_),
    .ZN(_3557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4024_ (.A1(_3543_),
    .A2(_3467_),
    .B(_3468_),
    .C(_3557_),
    .ZN(_3558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4025_ (.A1(_3452_),
    .A2(_3537_),
    .B(_3558_),
    .C(_3479_),
    .ZN(_3559_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4026_ (.A1(_3450_),
    .A2(_3529_),
    .B(_3559_),
    .C(_3484_),
    .ZN(_3560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4027_ (.A1(_3528_),
    .A2(_3313_),
    .B(_3315_),
    .C(_3560_),
    .ZN(_3561_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4028_ (.I(_3544_),
    .Z(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4029_ (.A1(_3368_),
    .A2(_3354_),
    .A3(_3562_),
    .ZN(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4030_ (.A1(_3297_),
    .A2(_3471_),
    .B(_3459_),
    .ZN(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4031_ (.I(_3446_),
    .Z(_3565_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4032_ (.A1(_3563_),
    .A2(_3564_),
    .B(_3565_),
    .ZN(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4033_ (.I(_3388_),
    .Z(_3567_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4034_ (.A1(_3545_),
    .A2(_3553_),
    .Z(_3568_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4035_ (.A1(_3388_),
    .A2(_3460_),
    .B(_3565_),
    .ZN(_3569_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4036_ (.A1(_3567_),
    .A2(_3568_),
    .B(_3569_),
    .ZN(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4037_ (.A1(_3566_),
    .A2(_3570_),
    .ZN(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4038_ (.A1(_3444_),
    .A2(_3571_),
    .B(_3488_),
    .ZN(_3572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4039_ (.A1(_3563_),
    .A2(_3564_),
    .B(_3489_),
    .ZN(_3573_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4040_ (.I(_3299_),
    .Z(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4041_ (.A1(_3299_),
    .A2(_3460_),
    .B(_3489_),
    .ZN(_3575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4042_ (.A1(_3574_),
    .A2(_3568_),
    .B(_3575_),
    .ZN(_3576_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4043_ (.A1(_3573_),
    .A2(_3576_),
    .Z(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4044_ (.A1(_3561_),
    .A2(_3572_),
    .B1(_3577_),
    .B2(_3443_),
    .ZN(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4045_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3562_),
    .Z(_3579_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4046_ (.A1(\as2650.holding_reg[2] ),
    .A2(_3562_),
    .ZN(_3580_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4047_ (.A1(_3579_),
    .A2(_3580_),
    .ZN(_3581_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4048_ (.I(_3581_),
    .Z(_3582_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4049_ (.A1(_3497_),
    .A2(_3445_),
    .ZN(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4050_ (.I(\as2650.psl[3] ),
    .ZN(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4051_ (.A1(_3584_),
    .A2(\as2650.carry ),
    .ZN(_3585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4052_ (.A1(_3421_),
    .A2(_3427_),
    .ZN(_3586_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4053_ (.A1(_3585_),
    .A2(_3402_),
    .B(_3586_),
    .ZN(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4054_ (.A1(_3500_),
    .A2(_3583_),
    .B1(_3508_),
    .B2(_3587_),
    .ZN(_3588_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4055_ (.A1(_3581_),
    .A2(_3588_),
    .Z(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4056_ (.A1(_3415_),
    .A2(_3589_),
    .ZN(_3590_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4057_ (.A1(_3497_),
    .A2(_3445_),
    .Z(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4058_ (.A1(_3591_),
    .A2(_3513_),
    .B(_3503_),
    .ZN(_3592_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _4059_ (.A1(_3581_),
    .A2(_3592_),
    .ZN(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4060_ (.I(\as2650.holding_reg[2] ),
    .Z(_0261_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4061_ (.I(_3257_),
    .Z(_0262_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4062_ (.I(_3458_),
    .Z(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4063_ (.A1(_3258_),
    .A2(_0263_),
    .ZN(_0264_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4064_ (.A1(_0261_),
    .A2(_0262_),
    .B(_0264_),
    .ZN(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4065_ (.A1(_3505_),
    .A2(_0265_),
    .ZN(_0266_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4066_ (.A1(_3407_),
    .A2(_3593_),
    .B(_0266_),
    .ZN(_0267_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4067_ (.A1(_3590_),
    .A2(_0267_),
    .B(_3164_),
    .ZN(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4068_ (.I(_3395_),
    .Z(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4069_ (.A1(_0261_),
    .A2(_3562_),
    .Z(_0270_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4070_ (.A1(_0269_),
    .A2(_3579_),
    .B(_0270_),
    .ZN(_0271_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4071_ (.A1(_3419_),
    .A2(_0271_),
    .B(_3397_),
    .ZN(_0272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4072_ (.A1(_3428_),
    .A2(_3582_),
    .B1(_0268_),
    .B2(_0272_),
    .ZN(_0273_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4073_ (.I(_0273_),
    .Z(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4074_ (.A1(_3436_),
    .A2(_0274_),
    .ZN(_0275_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4075_ (.A1(_3496_),
    .A2(_3578_),
    .B(_0275_),
    .ZN(_0276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4076_ (.A1(\as2650.r123[2][2] ),
    .A2(_3440_),
    .ZN(_0277_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4077_ (.A1(_3290_),
    .A2(_0276_),
    .B(_0277_),
    .ZN(_0002_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4078_ (.I(_3395_),
    .Z(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4079_ (.A1(_0278_),
    .A2(_3396_),
    .ZN(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4080_ (.A1(\as2650.holding_reg[3] ),
    .A2(_3535_),
    .ZN(_0280_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4081_ (.I(\as2650.holding_reg[3] ),
    .ZN(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4082_ (.A1(_3532_),
    .A2(_3534_),
    .Z(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4083_ (.I(_0282_),
    .Z(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4084_ (.A1(_0281_),
    .A2(_0283_),
    .ZN(_0284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4085_ (.A1(_0280_),
    .A2(_0284_),
    .ZN(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4086_ (.I(_0280_),
    .Z(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4087_ (.A1(_0286_),
    .A2(_0284_),
    .Z(_0287_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4088_ (.I(_0287_),
    .Z(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4089_ (.A1(_3591_),
    .A2(_3513_),
    .B(_3579_),
    .C(_3503_),
    .ZN(_0289_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4090_ (.A1(_3580_),
    .A2(_0289_),
    .ZN(_0290_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4091_ (.A1(_0288_),
    .A2(_0290_),
    .Z(_0291_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4092_ (.A1(_3408_),
    .A2(_0291_),
    .ZN(_0292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4093_ (.A1(_3499_),
    .A2(_3583_),
    .ZN(_0293_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4094_ (.A1(_3591_),
    .A2(_3509_),
    .B(_0293_),
    .ZN(_0294_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4095_ (.A1(_3581_),
    .A2(_0287_),
    .ZN(_0295_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4096_ (.A1(_0270_),
    .A2(_0265_),
    .A3(_0285_),
    .Z(_0296_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4097_ (.A1(_0294_),
    .A2(_0295_),
    .B(_0296_),
    .ZN(_0297_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4098_ (.A1(_0270_),
    .A2(_0265_),
    .ZN(_0298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4099_ (.A1(_3582_),
    .A2(_3588_),
    .B(_0288_),
    .C(_0298_),
    .ZN(_0299_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4100_ (.I(_3415_),
    .Z(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4101_ (.A1(_0297_),
    .A2(_0299_),
    .B(_0300_),
    .ZN(_0301_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4102_ (.A1(_0281_),
    .A2(_3261_),
    .ZN(_0302_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4103_ (.I(_3406_),
    .Z(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4104_ (.A1(_3261_),
    .A2(_3536_),
    .B(_0302_),
    .C(_0303_),
    .ZN(_0304_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4105_ (.I(_3404_),
    .Z(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4106_ (.I(_0282_),
    .Z(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4107_ (.A1(\as2650.holding_reg[3] ),
    .A2(_3258_),
    .ZN(_0307_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4108_ (.A1(_0262_),
    .A2(_0306_),
    .B(_0307_),
    .ZN(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4109_ (.A1(_0305_),
    .A2(_0308_),
    .ZN(_0309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4110_ (.I(_3164_),
    .Z(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__oai32_2 _4111_ (.A1(_0292_),
    .A2(_0301_),
    .A3(_0304_),
    .B1(_0309_),
    .B2(_0310_),
    .ZN(_0311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4112_ (.I(_3165_),
    .Z(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4113_ (.A1(_0312_),
    .A2(_0286_),
    .B(_3428_),
    .ZN(_0313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4114_ (.A1(_0311_),
    .A2(_0313_),
    .ZN(_0314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4115_ (.A1(_0279_),
    .A2(_0285_),
    .B(_0314_),
    .ZN(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4116_ (.I(_3300_),
    .Z(_0316_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4117_ (.I(_0306_),
    .Z(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4118_ (.A1(_3563_),
    .A2(_3536_),
    .Z(_0318_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4119_ (.I(_3298_),
    .Z(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4120_ (.A1(\as2650.idx_ctrl[1] ),
    .A2(_3186_),
    .ZN(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4121_ (.A1(_0263_),
    .A2(_3552_),
    .A3(_0283_),
    .Z(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4122_ (.A1(_3459_),
    .A2(_3553_),
    .B(_0306_),
    .ZN(_0322_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4123_ (.A1(_0320_),
    .A2(_0321_),
    .A3(_0322_),
    .ZN(_0323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4124_ (.A1(_0316_),
    .A2(_0317_),
    .B1(_0318_),
    .B2(_0319_),
    .C(_0323_),
    .ZN(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4125_ (.I(_0324_),
    .Z(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4126_ (.A1(_3310_),
    .A2(_0325_),
    .ZN(_0326_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _4127_ (.I(_3386_),
    .Z(_0327_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4128_ (.A1(_3385_),
    .A2(\as2650.addr_buff[6] ),
    .ZN(_0328_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4129_ (.A1(_0328_),
    .A2(_0321_),
    .A3(_0322_),
    .ZN(_0329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4130_ (.A1(_3389_),
    .A2(_0317_),
    .B1(_0318_),
    .B2(_0327_),
    .C(_0329_),
    .ZN(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4131_ (.I(_0330_),
    .Z(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4132_ (.I(_3546_),
    .Z(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4133_ (.I(_3323_),
    .Z(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__mux4_1 _4134_ (.I0(\as2650.r123[0][4] ),
    .I1(\as2650.r123[2][4] ),
    .I2(\as2650.r123_2[0][4] ),
    .I3(\as2650.r123_2[2][4] ),
    .S0(_3331_),
    .S1(_0333_),
    .Z(_0334_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4135_ (.A1(_3346_),
    .A2(_0334_),
    .ZN(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4136_ (.I(_3133_),
    .Z(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4137_ (.I0(\as2650.r123[1][4] ),
    .I1(\as2650.r123_2[1][4] ),
    .S(_3192_),
    .Z(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4138_ (.A1(\as2650.r0[4] ),
    .A2(_3197_),
    .Z(_0338_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4139_ (.A1(_0336_),
    .A2(_0337_),
    .B(_0338_),
    .C(_3135_),
    .ZN(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4140_ (.A1(_0335_),
    .A2(_0339_),
    .Z(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4141_ (.I(_0340_),
    .Z(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4142_ (.I(_0341_),
    .Z(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4143_ (.I(net4),
    .Z(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4144_ (.I(_0343_),
    .Z(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4145_ (.I(_0344_),
    .Z(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4146_ (.I(_0317_),
    .Z(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4147_ (.A1(_3281_),
    .A2(_3368_),
    .A3(_3354_),
    .A4(_3545_),
    .ZN(_0347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4148_ (.A1(_3545_),
    .A2(_3554_),
    .B(_0347_),
    .ZN(_0348_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4149_ (.A1(_0346_),
    .A2(_0348_),
    .Z(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4150_ (.A1(_3364_),
    .A2(_0349_),
    .ZN(_0350_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4151_ (.A1(_0345_),
    .A2(_3469_),
    .B(_3371_),
    .C(_0350_),
    .ZN(_0351_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4152_ (.A1(_3345_),
    .A2(_0342_),
    .B(_0351_),
    .C(_3377_),
    .ZN(_0352_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4153_ (.A1(_3318_),
    .A2(_0332_),
    .B(_0352_),
    .C(_3379_),
    .ZN(_0353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4154_ (.I(\as2650.r0[3] ),
    .Z(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4155_ (.I(_3276_),
    .Z(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4156_ (.I(_0355_),
    .Z(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4157_ (.I(_0356_),
    .Z(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4158_ (.A1(_3244_),
    .A2(_3250_),
    .ZN(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4159_ (.A1(_0357_),
    .A2(_3277_),
    .A3(_0358_),
    .ZN(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4160_ (.A1(_0354_),
    .A2(_0359_),
    .ZN(_0360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4161_ (.I(_3383_),
    .Z(_0361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4162_ (.A1(_0353_),
    .A2(_0360_),
    .B(_0361_),
    .ZN(_0362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4163_ (.A1(_3384_),
    .A2(_0331_),
    .B(_0362_),
    .C(_3442_),
    .ZN(_0363_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4164_ (.A1(_3436_),
    .A2(_0326_),
    .A3(_0363_),
    .ZN(_0364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4165_ (.A1(_3496_),
    .A2(_0315_),
    .B(_0364_),
    .ZN(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4166_ (.A1(\as2650.r123[2][3] ),
    .A2(_3440_),
    .ZN(_0366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4167_ (.A1(_3290_),
    .A2(_0365_),
    .B(_0366_),
    .ZN(_0003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4168_ (.I(_3289_),
    .Z(_0367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4169_ (.I(\as2650.holding_reg[4] ),
    .Z(_0368_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4170_ (.A1(_0335_),
    .A2(_0339_),
    .ZN(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4171_ (.I(_0369_),
    .Z(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4172_ (.A1(_0368_),
    .A2(_0370_),
    .ZN(_0371_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4173_ (.I(_0369_),
    .Z(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4174_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0372_),
    .Z(_0373_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4175_ (.A1(_0371_),
    .A2(_0373_),
    .Z(_0374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4176_ (.I(_0374_),
    .Z(_0375_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4177_ (.A1(_0286_),
    .A2(_0308_),
    .Z(_0376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_4 _4178_ (.A1(_0294_),
    .A2(_0295_),
    .B(_0376_),
    .C(_0296_),
    .ZN(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4179_ (.A1(_0374_),
    .A2(_0377_),
    .Z(_0378_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4180_ (.I(_3248_),
    .Z(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4181_ (.A1(_0368_),
    .A2(_0379_),
    .ZN(_0380_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4182_ (.A1(_0379_),
    .A2(_0341_),
    .B(_0380_),
    .C(_0300_),
    .ZN(_0381_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4183_ (.A1(_0300_),
    .A2(_0378_),
    .B(_0381_),
    .C(_3408_),
    .ZN(_0382_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4184_ (.I(_3512_),
    .Z(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4185_ (.I(_0284_),
    .ZN(_0384_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4186_ (.A1(_3580_),
    .A2(_0384_),
    .A3(_0289_),
    .B(_0286_),
    .ZN(_0385_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4187_ (.A1(_0374_),
    .A2(_0385_),
    .Z(_0386_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4188_ (.A1(\as2650.holding_reg[4] ),
    .A2(_0262_),
    .ZN(_0387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4189_ (.A1(_3246_),
    .A2(_0370_),
    .ZN(_0388_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4190_ (.A1(_0387_),
    .A2(_0388_),
    .Z(_0389_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4191_ (.A1(_0269_),
    .A2(_0389_),
    .ZN(_0390_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4192_ (.A1(_0383_),
    .A2(_0386_),
    .B1(_0390_),
    .B2(_3420_),
    .ZN(_0391_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4193_ (.A1(_0312_),
    .A2(_0371_),
    .B1(_0382_),
    .B2(_0391_),
    .ZN(_0392_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4194_ (.I0(_0375_),
    .I1(_0392_),
    .S(_0279_),
    .Z(_0393_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4195_ (.I(_0393_),
    .Z(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4196_ (.A1(_3296_),
    .A2(_3470_),
    .A3(_0263_),
    .A4(_0283_),
    .ZN(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4197_ (.I(_0395_),
    .Z(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4198_ (.A1(_0396_),
    .A2(_0341_),
    .Z(_0397_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4199_ (.A1(_0340_),
    .A2(_0321_),
    .Z(_0398_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _4200_ (.A1(_0319_),
    .A2(_0397_),
    .B1(_0398_),
    .B2(_3574_),
    .C1(_0316_),
    .C2(_0341_),
    .ZN(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4201_ (.I(_0399_),
    .Z(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4202_ (.A1(_3309_),
    .A2(_0400_),
    .ZN(_0401_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4203_ (.A1(_3565_),
    .A2(_0328_),
    .ZN(_0402_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4204_ (.I(_0370_),
    .Z(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4205_ (.A1(_0402_),
    .A2(_0403_),
    .ZN(_0404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4206_ (.A1(_0327_),
    .A2(_0397_),
    .B1(_0398_),
    .B2(_3567_),
    .C(_0404_),
    .ZN(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4207_ (.I(_0405_),
    .Z(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4208_ (.I0(\as2650.r123[2][5] ),
    .I1(\as2650.r123_2[2][5] ),
    .S(_3323_),
    .Z(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4209_ (.A1(_3136_),
    .A2(_0407_),
    .ZN(_0408_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4210_ (.A1(\as2650.r0[5] ),
    .A2(_3199_),
    .ZN(_0409_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4211_ (.I(\as2650.r123_2[0][5] ),
    .ZN(_0410_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4212_ (.A1(_3192_),
    .A2(_0410_),
    .ZN(_0411_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4213_ (.A1(_0333_),
    .A2(\as2650.r123[0][5] ),
    .B(_3333_),
    .C(_0411_),
    .ZN(_0412_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4214_ (.I(\as2650.r123_2[1][5] ),
    .ZN(_0413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4215_ (.A1(_3192_),
    .A2(_0413_),
    .ZN(_0414_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4216_ (.A1(_0333_),
    .A2(\as2650.r123[1][5] ),
    .B(_3326_),
    .C(_0414_),
    .ZN(_0415_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4217_ (.A1(_0408_),
    .A2(_0409_),
    .A3(_0412_),
    .A4(_0415_),
    .Z(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4218_ (.I(_0416_),
    .Z(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4219_ (.I(_0417_),
    .Z(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4220_ (.I(_0418_),
    .Z(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4221_ (.A1(_3549_),
    .A2(_3459_),
    .A3(_3553_),
    .A4(_0306_),
    .ZN(_0420_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4222_ (.A1(_0347_),
    .A2(_0317_),
    .B(_0420_),
    .ZN(_0421_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4223_ (.A1(_0403_),
    .A2(_0421_),
    .Z(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4224_ (.I(net5),
    .Z(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4225_ (.I(_0423_),
    .ZN(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4226_ (.I(_0424_),
    .Z(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4227_ (.A1(_0425_),
    .A2(_3365_),
    .ZN(_0426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4228_ (.A1(_3366_),
    .A2(_0422_),
    .B(_0426_),
    .C(_3371_),
    .ZN(_0427_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4229_ (.A1(_3345_),
    .A2(_0419_),
    .B(_0427_),
    .C(_3377_),
    .ZN(_0428_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4230_ (.A1(_3318_),
    .A2(_3537_),
    .B(_0428_),
    .C(_3379_),
    .ZN(_0429_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4231_ (.A1(\as2650.r0[4] ),
    .A2(_0359_),
    .ZN(_0430_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4232_ (.A1(_0429_),
    .A2(_0430_),
    .B(_0361_),
    .ZN(_0431_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4233_ (.A1(_3384_),
    .A2(_0406_),
    .B(_0431_),
    .C(_3442_),
    .ZN(_0432_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4234_ (.A1(_3436_),
    .A2(_0401_),
    .A3(_0432_),
    .ZN(_0433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4235_ (.A1(_3496_),
    .A2(_0394_),
    .B(_0433_),
    .ZN(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4236_ (.I(_3439_),
    .Z(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4237_ (.A1(\as2650.r123[2][4] ),
    .A2(_0435_),
    .ZN(_0436_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4238_ (.A1(_0367_),
    .A2(_0434_),
    .B(_0436_),
    .ZN(_0004_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4239_ (.I(_3494_),
    .Z(_0437_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4240_ (.I(_3428_),
    .Z(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4241_ (.A1(\as2650.holding_reg[5] ),
    .A2(_0416_),
    .Z(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4242_ (.A1(_0368_),
    .A2(_0403_),
    .Z(_0440_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4243_ (.A1(_0373_),
    .A2(_0385_),
    .B(_0440_),
    .ZN(_0441_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4244_ (.A1(_0439_),
    .A2(_0441_),
    .Z(_0442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4245_ (.A1(_0383_),
    .A2(_0442_),
    .ZN(_0443_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4246_ (.A1(_0278_),
    .A2(_3420_),
    .ZN(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4247_ (.A1(_0387_),
    .A2(_0388_),
    .ZN(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4248_ (.A1(_0371_),
    .A2(_0445_),
    .A3(_0439_),
    .ZN(_0446_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4249_ (.I(\as2650.holding_reg[5] ),
    .Z(_0447_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4250_ (.A1(_0408_),
    .A2(_0409_),
    .A3(_0412_),
    .A4(_0415_),
    .ZN(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4251_ (.I(_0448_),
    .Z(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4252_ (.A1(_0447_),
    .A2(_0449_),
    .Z(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4253_ (.A1(_0375_),
    .A2(_0377_),
    .A3(_0450_),
    .Z(_0451_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4254_ (.A1(_0375_),
    .A2(_0377_),
    .B1(_0389_),
    .B2(_0440_),
    .C(_0450_),
    .ZN(_0452_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _4255_ (.A1(_3506_),
    .A2(_0446_),
    .A3(_0451_),
    .A4(_0452_),
    .ZN(_0453_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4256_ (.A1(\as2650.holding_reg[5] ),
    .A2(_3246_),
    .Z(_0454_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4257_ (.A1(_3259_),
    .A2(_0449_),
    .B(_0454_),
    .ZN(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4258_ (.A1(_0303_),
    .A2(_0455_),
    .Z(_0456_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4259_ (.A1(_0444_),
    .A2(_0453_),
    .A3(_0456_),
    .Z(_0457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4260_ (.I(_0447_),
    .Z(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4261_ (.I(_0448_),
    .Z(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4262_ (.I(_0459_),
    .Z(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4263_ (.A1(_0458_),
    .A2(_0310_),
    .A3(_0460_),
    .ZN(_0461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4264_ (.A1(_0443_),
    .A2(_0457_),
    .B(_0461_),
    .C(_0312_),
    .ZN(_0462_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4265_ (.I(_0460_),
    .Z(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4266_ (.A1(_0458_),
    .A2(_0312_),
    .A3(_0463_),
    .Z(_0464_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4267_ (.A1(_0438_),
    .A2(_0439_),
    .ZN(_0465_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _4268_ (.A1(_0438_),
    .A2(_0462_),
    .A3(_0464_),
    .B(_0465_),
    .ZN(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4269_ (.I(_0466_),
    .ZN(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4270_ (.A1(_0395_),
    .A2(_0370_),
    .ZN(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4271_ (.A1(_0468_),
    .A2(_0449_),
    .Z(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4272_ (.A1(_0263_),
    .A2(_3552_),
    .A3(_0283_),
    .A4(_0340_),
    .ZN(_0470_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4273_ (.A1(_0470_),
    .A2(_0417_),
    .Z(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4274_ (.A1(_0320_),
    .A2(_0471_),
    .ZN(_0472_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4275_ (.A1(_3300_),
    .A2(_0418_),
    .Z(_0473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _4276_ (.A1(_0319_),
    .A2(_0469_),
    .B(_0472_),
    .C(_0473_),
    .ZN(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4277_ (.I(_0474_),
    .Z(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4278_ (.I(\as2650.r0[5] ),
    .Z(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4279_ (.I(_0372_),
    .Z(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4280_ (.A1(_3282_),
    .A2(_0396_),
    .A3(_0403_),
    .ZN(_0478_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4281_ (.A1(_0420_),
    .A2(_0477_),
    .B(_0478_),
    .ZN(_0479_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4282_ (.A1(_0460_),
    .A2(_0479_),
    .Z(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4283_ (.I(net6),
    .Z(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4284_ (.I(_0481_),
    .ZN(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4285_ (.I(_0482_),
    .Z(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4286_ (.A1(_0483_),
    .A2(_3469_),
    .B(_3371_),
    .ZN(_0484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4287_ (.A1(_3467_),
    .A2(_0480_),
    .B(_0484_),
    .ZN(_0485_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4288_ (.I0(\as2650.r123[2][6] ),
    .I1(\as2650.r123_2[2][6] ),
    .S(_0333_),
    .Z(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4289_ (.A1(_3137_),
    .A2(_0486_),
    .ZN(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4290_ (.A1(\as2650.r0[6] ),
    .A2(_3199_),
    .ZN(_0488_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4291_ (.I(\as2650.r123_2[0][6] ),
    .ZN(_0489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4292_ (.A1(_3324_),
    .A2(_0489_),
    .ZN(_0490_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4293_ (.A1(_3193_),
    .A2(\as2650.r123[0][6] ),
    .B(_3333_),
    .C(_0490_),
    .ZN(_0491_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4294_ (.I(\as2650.r123_2[1][6] ),
    .ZN(_0492_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4295_ (.A1(_3324_),
    .A2(_0492_),
    .ZN(_0493_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _4296_ (.A1(_3193_),
    .A2(\as2650.r123[1][6] ),
    .B(_3326_),
    .C(_0493_),
    .ZN(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4297_ (.A1(_0487_),
    .A2(_0488_),
    .A3(_0491_),
    .A4(_0494_),
    .ZN(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4298_ (.I(_0495_),
    .Z(_0496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4299_ (.I(_0496_),
    .Z(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4300_ (.A1(_3345_),
    .A2(_0497_),
    .B(_3377_),
    .ZN(_0498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4301_ (.A1(_0485_),
    .A2(_0498_),
    .ZN(_0499_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4302_ (.I(_0342_),
    .Z(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4303_ (.A1(_3479_),
    .A2(_0500_),
    .B(_3379_),
    .ZN(_0501_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4304_ (.A1(_0476_),
    .A2(_3484_),
    .B1(_0499_),
    .B2(_0501_),
    .C(_3315_),
    .ZN(_0502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4305_ (.A1(_0328_),
    .A2(_0471_),
    .ZN(_0503_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4306_ (.A1(_3389_),
    .A2(_0418_),
    .B1(_0469_),
    .B2(_0327_),
    .C(_0503_),
    .ZN(_0504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4307_ (.I(_0504_),
    .Z(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4308_ (.A1(_0361_),
    .A2(_0505_),
    .ZN(_0506_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4309_ (.A1(_3309_),
    .A2(_0502_),
    .A3(_0506_),
    .ZN(_0507_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4310_ (.A1(_3310_),
    .A2(_0475_),
    .B(_0507_),
    .ZN(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4311_ (.A1(_0437_),
    .A2(_0508_),
    .ZN(_0509_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4312_ (.A1(_0437_),
    .A2(_0467_),
    .B(_0509_),
    .ZN(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4313_ (.A1(\as2650.r123[2][5] ),
    .A2(_0435_),
    .ZN(_0511_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4314_ (.A1(_0367_),
    .A2(_0510_),
    .B(_0511_),
    .ZN(_0005_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4315_ (.A1(_0487_),
    .A2(_0488_),
    .A3(_0491_),
    .A4(_0494_),
    .Z(_0512_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4316_ (.A1(\as2650.holding_reg[6] ),
    .A2(_0512_),
    .Z(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4317_ (.I(_0513_),
    .Z(_0514_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4318_ (.A1(_0458_),
    .A2(_0460_),
    .ZN(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4319_ (.A1(_0447_),
    .A2(_0459_),
    .B1(_0373_),
    .B2(_0385_),
    .C(_0440_),
    .ZN(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4320_ (.A1(_0515_),
    .A2(_0516_),
    .ZN(_0517_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4321_ (.A1(_0514_),
    .A2(_0517_),
    .Z(_0518_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4322_ (.A1(_0447_),
    .A2(_0262_),
    .ZN(_0519_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4323_ (.A1(_3259_),
    .A2(_0417_),
    .B(_0519_),
    .ZN(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4324_ (.A1(_0455_),
    .A2(_0520_),
    .ZN(_0521_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4325_ (.A1(_0446_),
    .A2(_0521_),
    .Z(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4326_ (.A1(_0374_),
    .A2(_0377_),
    .A3(_0450_),
    .B(_0522_),
    .ZN(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4327_ (.A1(_0514_),
    .A2(_0523_),
    .Z(_0524_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4328_ (.I(_0512_),
    .Z(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4329_ (.A1(_3259_),
    .A2(_0525_),
    .ZN(_0526_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4330_ (.A1(\as2650.holding_reg[6] ),
    .A2(_3260_),
    .B(_0526_),
    .ZN(_0527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4331_ (.I(_0527_),
    .ZN(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _4332_ (.A1(_0300_),
    .A2(_0524_),
    .B1(_0528_),
    .B2(_0303_),
    .C(_0310_),
    .ZN(_0529_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4333_ (.A1(_0383_),
    .A2(_0518_),
    .B(_0529_),
    .ZN(_0530_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4334_ (.I(\as2650.holding_reg[6] ),
    .Z(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4335_ (.A1(_0531_),
    .A2(_0497_),
    .ZN(_0532_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4336_ (.A1(_0531_),
    .A2(_0497_),
    .B(_3517_),
    .ZN(_0533_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4337_ (.A1(_3423_),
    .A2(_0532_),
    .B(_0533_),
    .C(_0279_),
    .ZN(_0534_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4338_ (.A1(_0530_),
    .A2(_0534_),
    .ZN(_0535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4339_ (.A1(_0438_),
    .A2(_0514_),
    .B(_0535_),
    .ZN(_0536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4340_ (.I(_0536_),
    .Z(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4341_ (.A1(_0396_),
    .A2(_0372_),
    .A3(_0459_),
    .A4(_0496_),
    .ZN(_0538_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4342_ (.A1(_0468_),
    .A2(_0418_),
    .B(_0525_),
    .ZN(_0539_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4343_ (.A1(_0538_),
    .A2(_0539_),
    .ZN(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4344_ (.A1(_0340_),
    .A2(_0321_),
    .A3(_0417_),
    .ZN(_0541_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4345_ (.A1(_0541_),
    .A2(_0495_),
    .Z(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4346_ (.I(_0495_),
    .Z(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4347_ (.A1(_0402_),
    .A2(_0543_),
    .ZN(_0544_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4348_ (.A1(_0327_),
    .A2(_0540_),
    .B1(_0542_),
    .B2(_3567_),
    .C(_0544_),
    .ZN(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4349_ (.I(_0545_),
    .Z(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4350_ (.I(\as2650.r0[6] ),
    .Z(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4351_ (.A1(_0547_),
    .A2(_0359_),
    .ZN(_0548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4352_ (.I(_0463_),
    .Z(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4353_ (.I(_3340_),
    .Z(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4354_ (.A1(_3282_),
    .A2(_0396_),
    .A3(_0372_),
    .A4(_0449_),
    .Z(_0551_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4355_ (.A1(_0551_),
    .A2(_0543_),
    .ZN(_0552_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4356_ (.I(_0541_),
    .Z(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4357_ (.A1(_3473_),
    .A2(_0553_),
    .B1(_0538_),
    .B2(_3547_),
    .ZN(_0554_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4358_ (.A1(_3473_),
    .A2(_0553_),
    .A3(_0543_),
    .Z(_0555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _4359_ (.A1(_0552_),
    .A2(_0554_),
    .B(_0555_),
    .ZN(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4360_ (.I(net7),
    .Z(_0557_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4361_ (.I(_0557_),
    .ZN(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4362_ (.I(_0558_),
    .Z(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4363_ (.A1(_0559_),
    .A2(_3365_),
    .ZN(_0560_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4364_ (.A1(_3366_),
    .A2(_0556_),
    .B(_0560_),
    .C(_3468_),
    .ZN(_0561_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4365_ (.A1(_3452_),
    .A2(_0550_),
    .B(_0561_),
    .C(_3479_),
    .ZN(_0562_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4366_ (.A1(_3318_),
    .A2(_0549_),
    .B(_0562_),
    .C(_3484_),
    .ZN(_0563_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4367_ (.A1(_0548_),
    .A2(_0563_),
    .B(_3384_),
    .ZN(_0564_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4368_ (.A1(_3444_),
    .A2(_0546_),
    .B(_0564_),
    .ZN(_0565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4369_ (.I(_0525_),
    .Z(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4370_ (.A1(_3574_),
    .A2(_0542_),
    .Z(_0567_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _4371_ (.A1(_0316_),
    .A2(_0566_),
    .B1(_0540_),
    .B2(_0319_),
    .C(_0567_),
    .ZN(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4372_ (.I(_0568_),
    .Z(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4373_ (.A1(_3488_),
    .A2(_0569_),
    .ZN(_0570_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4374_ (.A1(_3443_),
    .A2(_0565_),
    .B(_0570_),
    .C(_3494_),
    .ZN(_0571_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4375_ (.A1(_0437_),
    .A2(_0537_),
    .B(_0571_),
    .ZN(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4376_ (.A1(\as2650.r123[2][6] ),
    .A2(_0435_),
    .ZN(_0573_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4377_ (.A1(_0367_),
    .A2(_0572_),
    .B(_0573_),
    .ZN(_0006_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4378_ (.A1(_3320_),
    .A2(_3322_),
    .A3(_3330_),
    .A4(_3336_),
    .ZN(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4379_ (.A1(\as2650.holding_reg[7] ),
    .A2(_0574_),
    .ZN(_0575_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4380_ (.I(\as2650.holding_reg[7] ),
    .ZN(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4381_ (.A1(_0576_),
    .A2(_3338_),
    .ZN(_0577_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4382_ (.A1(_0575_),
    .A2(_0577_),
    .ZN(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4383_ (.I(_0578_),
    .Z(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4384_ (.A1(_3247_),
    .A2(_0525_),
    .ZN(_0580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4385_ (.A1(_0531_),
    .A2(_3247_),
    .B(_0580_),
    .ZN(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4386_ (.A1(_0528_),
    .A2(_0581_),
    .ZN(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4387_ (.A1(_0513_),
    .A2(_0523_),
    .B(_0582_),
    .ZN(_0583_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4388_ (.A1(_0578_),
    .A2(_0583_),
    .Z(_0584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4389_ (.A1(_3261_),
    .A2(_0574_),
    .ZN(_0585_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4390_ (.A1(\as2650.holding_reg[7] ),
    .A2(_3248_),
    .ZN(_0586_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4391_ (.A1(_3415_),
    .A2(_0585_),
    .A3(_0586_),
    .Z(_0587_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4392_ (.A1(_3506_),
    .A2(_0584_),
    .B(_0587_),
    .C(_0383_),
    .ZN(_0588_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _4393_ (.A1(_0515_),
    .A2(_0513_),
    .A3(_0516_),
    .B(_0532_),
    .ZN(_0589_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4394_ (.A1(_0578_),
    .A2(_0589_),
    .Z(_0590_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4395_ (.A1(_3408_),
    .A2(_0590_),
    .B(_0444_),
    .ZN(_0591_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4396_ (.A1(_0576_),
    .A2(_3420_),
    .A3(_3340_),
    .ZN(_0592_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4397_ (.A1(_0588_),
    .A2(_0591_),
    .B(_0592_),
    .C(_3423_),
    .ZN(_0593_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4398_ (.A1(_3423_),
    .A2(_0575_),
    .ZN(_0594_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4399_ (.A1(_3398_),
    .A2(_0594_),
    .ZN(_0595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4400_ (.A1(_3398_),
    .A2(_0579_),
    .B1(_0593_),
    .B2(_0595_),
    .ZN(_0596_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4401_ (.I(_0596_),
    .Z(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4402_ (.A1(_0553_),
    .A2(_0496_),
    .ZN(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4403_ (.A1(_3338_),
    .A2(_0598_),
    .Z(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4404_ (.A1(_3337_),
    .A2(_0538_),
    .Z(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4405_ (.A1(_3565_),
    .A2(_0600_),
    .ZN(_0601_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4406_ (.A1(_3339_),
    .A2(_3389_),
    .B1(_0599_),
    .B2(_3567_),
    .C(_0601_),
    .ZN(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4407_ (.I(_0602_),
    .Z(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4408_ (.I(_0566_),
    .Z(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _4409_ (.A1(_3473_),
    .A2(_0470_),
    .A3(_0459_),
    .A4(_0496_),
    .ZN(_0605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4410_ (.A1(_0551_),
    .A2(_0543_),
    .B(_0605_),
    .ZN(_0606_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_2 _4411_ (.A1(_3338_),
    .A2(_0606_),
    .Z(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4412_ (.A1(_3366_),
    .A2(_0607_),
    .ZN(_0608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4413_ (.I(net8),
    .Z(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4414_ (.I(_0609_),
    .Z(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4415_ (.I(_0610_),
    .Z(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4416_ (.A1(_0611_),
    .A2(_3467_),
    .B(_3468_),
    .ZN(_0612_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4417_ (.A1(_3584_),
    .A2(_3369_),
    .B(_3403_),
    .ZN(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _4418_ (.A1(_0608_),
    .A2(_0612_),
    .B1(_0613_),
    .B2(_3452_),
    .ZN(_0614_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4419_ (.A1(_3450_),
    .A2(_0614_),
    .ZN(_0615_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4420_ (.A1(_3450_),
    .A2(_0604_),
    .B(_0615_),
    .C(_3313_),
    .ZN(_0616_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4421_ (.I(\as2650.r0[7] ),
    .Z(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4422_ (.I(_0617_),
    .ZN(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4423_ (.A1(_0618_),
    .A2(_0359_),
    .B(_0361_),
    .ZN(_0619_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4424_ (.A1(_3444_),
    .A2(_0603_),
    .B1(_0616_),
    .B2(_0619_),
    .ZN(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4425_ (.A1(_3489_),
    .A2(_0600_),
    .ZN(_0621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _4426_ (.A1(_3339_),
    .A2(_0316_),
    .B1(_0599_),
    .B2(_3574_),
    .C(_0621_),
    .ZN(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4427_ (.I(_0622_),
    .Z(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4428_ (.A1(_3488_),
    .A2(_0623_),
    .ZN(_0624_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4429_ (.A1(_3443_),
    .A2(_0620_),
    .B(_0624_),
    .C(_3494_),
    .ZN(_0625_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4430_ (.A1(_0437_),
    .A2(_0597_),
    .B(_0625_),
    .ZN(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4431_ (.A1(\as2650.r123[2][7] ),
    .A2(_0435_),
    .ZN(_0627_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4432_ (.A1(_0367_),
    .A2(_0626_),
    .B(_0627_),
    .ZN(_0007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4433_ (.A1(_3288_),
    .A2(_3327_),
    .ZN(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4434_ (.I(_0628_),
    .Z(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4435_ (.A1(_3288_),
    .A2(_3327_),
    .B(_3438_),
    .ZN(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4436_ (.I(_0630_),
    .Z(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4437_ (.A1(\as2650.r123[1][0] ),
    .A2(_0631_),
    .ZN(_0632_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4438_ (.A1(_3437_),
    .A2(_0629_),
    .B(_0632_),
    .ZN(_0008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4439_ (.A1(\as2650.r123[1][1] ),
    .A2(_0631_),
    .ZN(_0633_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4440_ (.A1(_3526_),
    .A2(_0629_),
    .B(_0633_),
    .ZN(_0009_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4441_ (.A1(\as2650.r123[1][2] ),
    .A2(_0631_),
    .ZN(_0634_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4442_ (.A1(_0276_),
    .A2(_0629_),
    .B(_0634_),
    .ZN(_0010_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4443_ (.A1(\as2650.r123[1][3] ),
    .A2(_0631_),
    .ZN(_0635_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4444_ (.A1(_0365_),
    .A2(_0629_),
    .B(_0635_),
    .ZN(_0011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4445_ (.I(_0628_),
    .Z(_0636_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4446_ (.I(_0630_),
    .Z(_0637_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4447_ (.A1(\as2650.r123[1][4] ),
    .A2(_0637_),
    .ZN(_0638_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4448_ (.A1(_0434_),
    .A2(_0636_),
    .B(_0638_),
    .ZN(_0012_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4449_ (.A1(\as2650.r123[1][5] ),
    .A2(_0637_),
    .ZN(_0639_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4450_ (.A1(_0510_),
    .A2(_0636_),
    .B(_0639_),
    .ZN(_0013_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4451_ (.A1(\as2650.r123[1][6] ),
    .A2(_0637_),
    .ZN(_0640_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4452_ (.A1(_0572_),
    .A2(_0636_),
    .B(_0640_),
    .ZN(_0014_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4453_ (.A1(\as2650.r123[1][7] ),
    .A2(_0637_),
    .ZN(_0641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4454_ (.A1(_0626_),
    .A2(_0636_),
    .B(_0641_),
    .ZN(_0015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4455_ (.I(\as2650.pc[0] ),
    .Z(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4456_ (.I(_0642_),
    .Z(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4457_ (.I(_0643_),
    .ZN(_0644_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4458_ (.I(_0644_),
    .Z(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4459_ (.I(_0645_),
    .Z(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4460_ (.I(_0646_),
    .Z(_0647_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4461_ (.A1(\as2650.stack_ptr[1] ),
    .A2(\as2650.stack_ptr[0] ),
    .ZN(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4462_ (.I(_0648_),
    .Z(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4463_ (.I(_0649_),
    .Z(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4464_ (.I(_0650_),
    .Z(_0651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4465_ (.I(\as2650.stack_ptr[2] ),
    .Z(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4466_ (.I(_3140_),
    .Z(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4467_ (.A1(_3206_),
    .A2(_3361_),
    .ZN(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4468_ (.I(_3216_),
    .ZN(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4469_ (.A1(_3215_),
    .A2(_0655_),
    .A3(_3213_),
    .ZN(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4470_ (.A1(_3304_),
    .A2(_0656_),
    .ZN(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4471_ (.I(\as2650.addr_buff[7] ),
    .Z(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4472_ (.I(_0658_),
    .Z(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4473_ (.I(_3181_),
    .Z(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4474_ (.I(_3180_),
    .Z(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4475_ (.A1(_3268_),
    .A2(_3217_),
    .A3(_0661_),
    .A4(_3214_),
    .ZN(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4476_ (.A1(_0660_),
    .A2(_0662_),
    .Z(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4477_ (.I(_0663_),
    .Z(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4478_ (.A1(_0659_),
    .A2(_0664_),
    .ZN(_0665_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4479_ (.A1(_0654_),
    .A2(_0657_),
    .A3(_0665_),
    .ZN(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4480_ (.A1(_3256_),
    .A2(_0278_),
    .A3(_3242_),
    .ZN(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4481_ (.I(_3279_),
    .Z(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4482_ (.I(_0668_),
    .Z(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4483_ (.A1(_3202_),
    .A2(_3178_),
    .ZN(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4484_ (.A1(_3138_),
    .A2(_3405_),
    .A3(_0670_),
    .ZN(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4485_ (.I(_0671_),
    .Z(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4486_ (.I(_0672_),
    .Z(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4487_ (.A1(_0669_),
    .A2(_0673_),
    .ZN(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4488_ (.I(_3206_),
    .Z(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4489_ (.I(_3197_),
    .Z(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4490_ (.I(_3346_),
    .Z(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4491_ (.A1(_0676_),
    .A2(_0677_),
    .ZN(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4492_ (.A1(_3154_),
    .A2(_3171_),
    .ZN(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4493_ (.A1(_0678_),
    .A2(_3505_),
    .A3(_0679_),
    .ZN(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4494_ (.A1(_0675_),
    .A2(_0680_),
    .ZN(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4495_ (.I(_0681_),
    .Z(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4496_ (.I(_0661_),
    .Z(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4497_ (.A1(_3267_),
    .A2(_3216_),
    .A3(_3213_),
    .Z(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4498_ (.I(_0684_),
    .Z(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4499_ (.A1(_0683_),
    .A2(_3274_),
    .A3(_0685_),
    .ZN(_0686_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4500_ (.I(_0686_),
    .Z(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__oai33_1 _4501_ (.A1(_0666_),
    .A2(_0667_),
    .A3(_0674_),
    .B1(_0682_),
    .B2(_0305_),
    .B3(_0687_),
    .ZN(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4502_ (.A1(_0652_),
    .A2(_0653_),
    .A3(_0688_),
    .Z(_0689_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4503_ (.A1(_0651_),
    .A2(_0689_),
    .ZN(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4504_ (.I(_0690_),
    .Z(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4505_ (.I(_0691_),
    .Z(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4506_ (.I(_0690_),
    .Z(_0693_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4507_ (.A1(\as2650.stack[4][0] ),
    .A2(_0693_),
    .ZN(_0694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4508_ (.A1(_0647_),
    .A2(_0692_),
    .B(_0694_),
    .ZN(_0016_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4509_ (.I(\as2650.pc[1] ),
    .ZN(_0695_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4510_ (.I(_0695_),
    .Z(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4511_ (.I(_0696_),
    .Z(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4512_ (.A1(\as2650.stack[4][1] ),
    .A2(_0693_),
    .ZN(_0698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4513_ (.A1(_0697_),
    .A2(_0692_),
    .B(_0698_),
    .ZN(_0017_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4514_ (.I(\as2650.pc[2] ),
    .ZN(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4515_ (.I(_0699_),
    .Z(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4516_ (.I(_0700_),
    .Z(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4517_ (.I(_0701_),
    .Z(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4518_ (.A1(\as2650.stack[4][2] ),
    .A2(_0693_),
    .ZN(_0703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4519_ (.A1(_0702_),
    .A2(_0692_),
    .B(_0703_),
    .ZN(_0018_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _4520_ (.I(\as2650.pc[3] ),
    .ZN(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4521_ (.I(_0704_),
    .Z(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4522_ (.I(_0705_),
    .Z(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4523_ (.A1(\as2650.stack[4][3] ),
    .A2(_0693_),
    .ZN(_0707_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4524_ (.A1(_0706_),
    .A2(_0692_),
    .B(_0707_),
    .ZN(_0019_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4525_ (.I(\as2650.pc[4] ),
    .ZN(_0708_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4526_ (.I(_0708_),
    .Z(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4527_ (.I(_0709_),
    .Z(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4528_ (.I(_0710_),
    .Z(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4529_ (.I(_0691_),
    .Z(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4530_ (.I(_0690_),
    .Z(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4531_ (.A1(\as2650.stack[4][4] ),
    .A2(_0713_),
    .ZN(_0714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4532_ (.A1(_0711_),
    .A2(_0712_),
    .B(_0714_),
    .ZN(_0020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4533_ (.I(\as2650.pc[5] ),
    .Z(_0715_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4534_ (.I(_0715_),
    .ZN(_0716_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4535_ (.I(_0716_),
    .Z(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4536_ (.I(_0717_),
    .Z(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4537_ (.A1(\as2650.stack[4][5] ),
    .A2(_0713_),
    .ZN(_0719_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4538_ (.A1(_0718_),
    .A2(_0712_),
    .B(_0719_),
    .ZN(_0021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4539_ (.I(\as2650.pc[6] ),
    .Z(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4540_ (.I(_0720_),
    .ZN(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4541_ (.I(_0721_),
    .Z(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4542_ (.A1(\as2650.stack[4][6] ),
    .A2(_0713_),
    .ZN(_0723_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4543_ (.A1(_0722_),
    .A2(_0712_),
    .B(_0723_),
    .ZN(_0022_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4544_ (.I(\as2650.pc[7] ),
    .ZN(_0724_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4545_ (.I(_0724_),
    .Z(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4546_ (.I(_0725_),
    .Z(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4547_ (.A1(\as2650.stack[4][7] ),
    .A2(_0713_),
    .ZN(_0727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4548_ (.A1(_0726_),
    .A2(_0712_),
    .B(_0727_),
    .ZN(_0023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4549_ (.I(\as2650.pc[8] ),
    .Z(_0728_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4550_ (.I(_0728_),
    .Z(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4551_ (.I(_0729_),
    .Z(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4552_ (.I(_0730_),
    .Z(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4553_ (.I0(_0731_),
    .I1(\as2650.stack[4][8] ),
    .S(_0691_),
    .Z(_0732_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4554_ (.I(_0732_),
    .Z(_0024_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4555_ (.I(\as2650.pc[9] ),
    .ZN(_0733_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4556_ (.I(_0733_),
    .Z(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4557_ (.I(_0734_),
    .Z(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4558_ (.I(_0691_),
    .Z(_0736_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4559_ (.I(_0690_),
    .Z(_0737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4560_ (.A1(\as2650.stack[4][9] ),
    .A2(_0737_),
    .ZN(_0738_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4561_ (.A1(_0735_),
    .A2(_0736_),
    .B(_0738_),
    .ZN(_0025_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4562_ (.I(\as2650.pc[10] ),
    .ZN(_0739_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4563_ (.I(_0739_),
    .Z(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4564_ (.I(_0740_),
    .Z(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4565_ (.A1(\as2650.stack[4][10] ),
    .A2(_0737_),
    .ZN(_0742_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4566_ (.A1(_0741_),
    .A2(_0736_),
    .B(_0742_),
    .ZN(_0026_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4567_ (.I(\as2650.pc[11] ),
    .ZN(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4568_ (.I(_0743_),
    .Z(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4569_ (.I(_0744_),
    .Z(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4570_ (.A1(\as2650.stack[4][11] ),
    .A2(_0737_),
    .ZN(_0746_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4571_ (.A1(_0745_),
    .A2(_0736_),
    .B(_0746_),
    .ZN(_0027_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4572_ (.I(\as2650.pc[12] ),
    .ZN(_0747_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4573_ (.I(_0747_),
    .Z(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4574_ (.I(_0748_),
    .Z(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4575_ (.A1(\as2650.stack[4][12] ),
    .A2(_0737_),
    .ZN(_0750_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4576_ (.A1(_0749_),
    .A2(_0736_),
    .B(_0750_),
    .ZN(_0028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4577_ (.I(\as2650.stack_ptr[0] ),
    .Z(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4578_ (.A1(\as2650.stack_ptr[1] ),
    .A2(_0751_),
    .Z(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4579_ (.I(_0752_),
    .Z(_0753_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4580_ (.I(_0753_),
    .Z(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4581_ (.I(_0754_),
    .Z(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4582_ (.A1(_0653_),
    .A2(_0688_),
    .ZN(_0756_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4583_ (.A1(_0652_),
    .A2(_0756_),
    .ZN(_0757_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4584_ (.A1(_0755_),
    .A2(_0757_),
    .ZN(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4585_ (.I(_0758_),
    .Z(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4586_ (.I(_0759_),
    .Z(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4587_ (.I(_0758_),
    .Z(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4588_ (.A1(\as2650.stack[3][0] ),
    .A2(_0761_),
    .ZN(_0762_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4589_ (.A1(_0647_),
    .A2(_0760_),
    .B(_0762_),
    .ZN(_0029_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4590_ (.A1(\as2650.stack[3][1] ),
    .A2(_0761_),
    .ZN(_0763_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4591_ (.A1(_0697_),
    .A2(_0760_),
    .B(_0763_),
    .ZN(_0030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4592_ (.A1(\as2650.stack[3][2] ),
    .A2(_0761_),
    .ZN(_0764_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4593_ (.A1(_0702_),
    .A2(_0760_),
    .B(_0764_),
    .ZN(_0031_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4594_ (.A1(\as2650.stack[3][3] ),
    .A2(_0761_),
    .ZN(_0765_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4595_ (.A1(_0706_),
    .A2(_0760_),
    .B(_0765_),
    .ZN(_0032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4596_ (.I(_0759_),
    .Z(_0766_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4597_ (.I(_0758_),
    .Z(_0767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4598_ (.A1(\as2650.stack[3][4] ),
    .A2(_0767_),
    .ZN(_0768_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4599_ (.A1(_0711_),
    .A2(_0766_),
    .B(_0768_),
    .ZN(_0033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4600_ (.A1(\as2650.stack[3][5] ),
    .A2(_0767_),
    .ZN(_0769_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4601_ (.A1(_0718_),
    .A2(_0766_),
    .B(_0769_),
    .ZN(_0034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4602_ (.A1(\as2650.stack[3][6] ),
    .A2(_0767_),
    .ZN(_0770_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4603_ (.A1(_0722_),
    .A2(_0766_),
    .B(_0770_),
    .ZN(_0035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4604_ (.A1(\as2650.stack[3][7] ),
    .A2(_0767_),
    .ZN(_0771_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4605_ (.A1(_0726_),
    .A2(_0766_),
    .B(_0771_),
    .ZN(_0036_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4606_ (.I0(_0731_),
    .I1(\as2650.stack[3][8] ),
    .S(_0759_),
    .Z(_0772_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4607_ (.I(_0772_),
    .Z(_0037_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4608_ (.I(_0759_),
    .Z(_0773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4609_ (.I(_0758_),
    .Z(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4610_ (.A1(\as2650.stack[3][9] ),
    .A2(_0774_),
    .ZN(_0775_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4611_ (.A1(_0735_),
    .A2(_0773_),
    .B(_0775_),
    .ZN(_0038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4612_ (.A1(\as2650.stack[3][10] ),
    .A2(_0774_),
    .ZN(_0776_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4613_ (.A1(_0741_),
    .A2(_0773_),
    .B(_0776_),
    .ZN(_0039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4614_ (.A1(\as2650.stack[3][11] ),
    .A2(_0774_),
    .ZN(_0777_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4615_ (.A1(_0745_),
    .A2(_0773_),
    .B(_0777_),
    .ZN(_0040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4616_ (.A1(\as2650.stack[3][12] ),
    .A2(_0774_),
    .ZN(_0778_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4617_ (.A1(_0749_),
    .A2(_0773_),
    .B(_0778_),
    .ZN(_0041_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4618_ (.I(\as2650.stack_ptr[1] ),
    .ZN(_0779_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4619_ (.A1(_0779_),
    .A2(_0751_),
    .ZN(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4620_ (.I(_0780_),
    .Z(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4621_ (.I(_0781_),
    .Z(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4622_ (.A1(_0757_),
    .A2(_0782_),
    .ZN(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4623_ (.I(_0783_),
    .Z(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4624_ (.I(_0784_),
    .Z(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4625_ (.I(_0783_),
    .Z(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4626_ (.A1(\as2650.stack[2][0] ),
    .A2(_0786_),
    .ZN(_0787_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4627_ (.A1(_0647_),
    .A2(_0785_),
    .B(_0787_),
    .ZN(_0042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4628_ (.A1(\as2650.stack[2][1] ),
    .A2(_0786_),
    .ZN(_0788_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4629_ (.A1(_0697_),
    .A2(_0785_),
    .B(_0788_),
    .ZN(_0043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4630_ (.A1(\as2650.stack[2][2] ),
    .A2(_0786_),
    .ZN(_0789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4631_ (.A1(_0702_),
    .A2(_0785_),
    .B(_0789_),
    .ZN(_0044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4632_ (.A1(\as2650.stack[2][3] ),
    .A2(_0786_),
    .ZN(_0790_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4633_ (.A1(_0706_),
    .A2(_0785_),
    .B(_0790_),
    .ZN(_0045_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4634_ (.I(_0784_),
    .Z(_0791_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4635_ (.I(_0783_),
    .Z(_0792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4636_ (.A1(\as2650.stack[2][4] ),
    .A2(_0792_),
    .ZN(_0793_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4637_ (.A1(_0711_),
    .A2(_0791_),
    .B(_0793_),
    .ZN(_0046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4638_ (.A1(\as2650.stack[2][5] ),
    .A2(_0792_),
    .ZN(_0794_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4639_ (.A1(_0718_),
    .A2(_0791_),
    .B(_0794_),
    .ZN(_0047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4640_ (.A1(\as2650.stack[2][6] ),
    .A2(_0792_),
    .ZN(_0795_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4641_ (.A1(_0722_),
    .A2(_0791_),
    .B(_0795_),
    .ZN(_0048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4642_ (.A1(\as2650.stack[2][7] ),
    .A2(_0792_),
    .ZN(_0796_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4643_ (.A1(_0726_),
    .A2(_0791_),
    .B(_0796_),
    .ZN(_0049_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4644_ (.I0(_0731_),
    .I1(\as2650.stack[2][8] ),
    .S(_0784_),
    .Z(_0797_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4645_ (.I(_0797_),
    .Z(_0050_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4646_ (.I(_0784_),
    .Z(_0798_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4647_ (.I(_0783_),
    .Z(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4648_ (.A1(\as2650.stack[2][9] ),
    .A2(_0799_),
    .ZN(_0800_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4649_ (.A1(_0735_),
    .A2(_0798_),
    .B(_0800_),
    .ZN(_0051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4650_ (.A1(\as2650.stack[2][10] ),
    .A2(_0799_),
    .ZN(_0801_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4651_ (.A1(_0741_),
    .A2(_0798_),
    .B(_0801_),
    .ZN(_0052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4652_ (.A1(\as2650.stack[2][11] ),
    .A2(_0799_),
    .ZN(_0802_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4653_ (.A1(_0745_),
    .A2(_0798_),
    .B(_0802_),
    .ZN(_0053_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4654_ (.A1(\as2650.stack[2][12] ),
    .A2(_0799_),
    .ZN(_0803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4655_ (.A1(_0749_),
    .A2(_0798_),
    .B(_0803_),
    .ZN(_0054_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4656_ (.A1(_0779_),
    .A2(\as2650.stack_ptr[0] ),
    .Z(_0804_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4657_ (.I(_0804_),
    .Z(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4658_ (.I(_0805_),
    .Z(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4659_ (.A1(_0757_),
    .A2(_0806_),
    .ZN(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4660_ (.I(_0807_),
    .Z(_0808_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4661_ (.I(_0808_),
    .Z(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4662_ (.I(_0807_),
    .Z(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4663_ (.A1(\as2650.stack[1][0] ),
    .A2(_0810_),
    .ZN(_0811_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4664_ (.A1(_0647_),
    .A2(_0809_),
    .B(_0811_),
    .ZN(_0055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4665_ (.A1(\as2650.stack[1][1] ),
    .A2(_0810_),
    .ZN(_0812_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4666_ (.A1(_0697_),
    .A2(_0809_),
    .B(_0812_),
    .ZN(_0056_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4667_ (.I(_0701_),
    .Z(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4668_ (.A1(\as2650.stack[1][2] ),
    .A2(_0810_),
    .ZN(_0814_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4669_ (.A1(_0813_),
    .A2(_0809_),
    .B(_0814_),
    .ZN(_0057_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4670_ (.I(_0705_),
    .Z(_0815_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4671_ (.A1(\as2650.stack[1][3] ),
    .A2(_0810_),
    .ZN(_0816_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4672_ (.A1(_0815_),
    .A2(_0809_),
    .B(_0816_),
    .ZN(_0058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4673_ (.I(_0710_),
    .Z(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4674_ (.I(_0808_),
    .Z(_0818_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4675_ (.I(_0807_),
    .Z(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4676_ (.A1(\as2650.stack[1][4] ),
    .A2(_0819_),
    .ZN(_0820_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4677_ (.A1(_0817_),
    .A2(_0818_),
    .B(_0820_),
    .ZN(_0059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4678_ (.I(_0717_),
    .Z(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4679_ (.A1(\as2650.stack[1][5] ),
    .A2(_0819_),
    .ZN(_0822_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4680_ (.A1(_0821_),
    .A2(_0818_),
    .B(_0822_),
    .ZN(_0060_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4681_ (.I(_0721_),
    .Z(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4682_ (.A1(\as2650.stack[1][6] ),
    .A2(_0819_),
    .ZN(_0824_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4683_ (.A1(_0823_),
    .A2(_0818_),
    .B(_0824_),
    .ZN(_0061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4684_ (.A1(\as2650.stack[1][7] ),
    .A2(_0819_),
    .ZN(_0825_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4685_ (.A1(_0726_),
    .A2(_0818_),
    .B(_0825_),
    .ZN(_0062_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4686_ (.I0(_0731_),
    .I1(\as2650.stack[1][8] ),
    .S(_0808_),
    .Z(_0826_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4687_ (.I(_0826_),
    .Z(_0063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4688_ (.I(_0734_),
    .Z(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4689_ (.I(_0808_),
    .Z(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4690_ (.I(_0807_),
    .Z(_0829_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4691_ (.A1(\as2650.stack[1][9] ),
    .A2(_0829_),
    .ZN(_0830_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4692_ (.A1(_0827_),
    .A2(_0828_),
    .B(_0830_),
    .ZN(_0064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4693_ (.I(_0740_),
    .Z(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4694_ (.A1(\as2650.stack[1][10] ),
    .A2(_0829_),
    .ZN(_0832_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4695_ (.A1(_0831_),
    .A2(_0828_),
    .B(_0832_),
    .ZN(_0065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4696_ (.A1(\as2650.stack[1][11] ),
    .A2(_0829_),
    .ZN(_0833_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4697_ (.A1(_0745_),
    .A2(_0828_),
    .B(_0833_),
    .ZN(_0066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4698_ (.A1(\as2650.stack[1][12] ),
    .A2(_0829_),
    .ZN(_0834_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4699_ (.A1(_0749_),
    .A2(_0828_),
    .B(_0834_),
    .ZN(_0067_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4700_ (.I(_0646_),
    .Z(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4701_ (.A1(_0651_),
    .A2(_0757_),
    .ZN(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4702_ (.I(_0836_),
    .Z(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4703_ (.I(_0837_),
    .Z(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4704_ (.I(_0836_),
    .Z(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4705_ (.A1(\as2650.stack[0][0] ),
    .A2(_0839_),
    .ZN(_0840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4706_ (.A1(_0835_),
    .A2(_0838_),
    .B(_0840_),
    .ZN(_0068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4707_ (.I(_0696_),
    .Z(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4708_ (.A1(\as2650.stack[0][1] ),
    .A2(_0839_),
    .ZN(_0842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4709_ (.A1(_0841_),
    .A2(_0838_),
    .B(_0842_),
    .ZN(_0069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4710_ (.A1(\as2650.stack[0][2] ),
    .A2(_0839_),
    .ZN(_0843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4711_ (.A1(_0813_),
    .A2(_0838_),
    .B(_0843_),
    .ZN(_0070_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4712_ (.A1(\as2650.stack[0][3] ),
    .A2(_0839_),
    .ZN(_0844_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4713_ (.A1(_0815_),
    .A2(_0838_),
    .B(_0844_),
    .ZN(_0071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4714_ (.I(_0837_),
    .Z(_0845_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4715_ (.I(_0836_),
    .Z(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4716_ (.A1(\as2650.stack[0][4] ),
    .A2(_0846_),
    .ZN(_0847_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4717_ (.A1(_0817_),
    .A2(_0845_),
    .B(_0847_),
    .ZN(_0072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4718_ (.A1(\as2650.stack[0][5] ),
    .A2(_0846_),
    .ZN(_0848_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4719_ (.A1(_0821_),
    .A2(_0845_),
    .B(_0848_),
    .ZN(_0073_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4720_ (.A1(\as2650.stack[0][6] ),
    .A2(_0846_),
    .ZN(_0849_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4721_ (.A1(_0823_),
    .A2(_0845_),
    .B(_0849_),
    .ZN(_0074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4722_ (.I(_0725_),
    .Z(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4723_ (.A1(\as2650.stack[0][7] ),
    .A2(_0846_),
    .ZN(_0851_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4724_ (.A1(_0850_),
    .A2(_0845_),
    .B(_0851_),
    .ZN(_0075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4725_ (.I(_0730_),
    .Z(_0852_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4726_ (.I0(_0852_),
    .I1(\as2650.stack[0][8] ),
    .S(_0837_),
    .Z(_0853_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4727_ (.I(_0853_),
    .Z(_0076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4728_ (.I(_0837_),
    .Z(_0854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4729_ (.I(_0836_),
    .Z(_0855_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4730_ (.A1(\as2650.stack[0][9] ),
    .A2(_0855_),
    .ZN(_0856_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4731_ (.A1(_0827_),
    .A2(_0854_),
    .B(_0856_),
    .ZN(_0077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4732_ (.A1(\as2650.stack[0][10] ),
    .A2(_0855_),
    .ZN(_0857_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4733_ (.A1(_0831_),
    .A2(_0854_),
    .B(_0857_),
    .ZN(_0078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4734_ (.I(_0744_),
    .Z(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4735_ (.A1(\as2650.stack[0][11] ),
    .A2(_0855_),
    .ZN(_0859_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4736_ (.A1(_0858_),
    .A2(_0854_),
    .B(_0859_),
    .ZN(_0079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4737_ (.I(_0748_),
    .Z(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4738_ (.A1(\as2650.stack[0][12] ),
    .A2(_0855_),
    .ZN(_0861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4739_ (.A1(_0860_),
    .A2(_0854_),
    .B(_0861_),
    .ZN(_0080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4740_ (.I(_3254_),
    .Z(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4741_ (.I(_0862_),
    .Z(_0863_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4742_ (.I(_0863_),
    .Z(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4743_ (.A1(_3195_),
    .A2(_3139_),
    .ZN(_0865_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4744_ (.A1(_0864_),
    .A2(_3272_),
    .A3(_0865_),
    .ZN(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4745_ (.I(_0866_),
    .Z(_0867_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4746_ (.I(_3135_),
    .Z(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4747_ (.A1(_0336_),
    .A2(_0868_),
    .ZN(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4748_ (.A1(_3253_),
    .A2(_0869_),
    .A3(_3139_),
    .ZN(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4749_ (.I(_0870_),
    .Z(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4750_ (.A1(_3188_),
    .A2(_0871_),
    .ZN(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4751_ (.I(_0872_),
    .Z(_0873_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4752_ (.A1(_3200_),
    .A2(_0865_),
    .ZN(_0874_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4753_ (.I(_0874_),
    .Z(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4754_ (.A1(_3227_),
    .A2(_3232_),
    .A3(_0875_),
    .ZN(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4755_ (.I(_0876_),
    .Z(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4756_ (.I(_0877_),
    .Z(_0878_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4757_ (.I(_3374_),
    .Z(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4758_ (.A1(_3208_),
    .A2(_3211_),
    .ZN(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4759_ (.A1(_0880_),
    .A2(_0654_),
    .ZN(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4760_ (.A1(_3279_),
    .A2(_0881_),
    .A3(_0870_),
    .ZN(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4761_ (.I(_0882_),
    .Z(_0883_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4762_ (.I(_3358_),
    .Z(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4763_ (.A1(_3214_),
    .A2(_3220_),
    .ZN(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4764_ (.A1(_3169_),
    .A2(_0884_),
    .A3(_0885_),
    .A4(_0870_),
    .ZN(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4765_ (.A1(_3175_),
    .A2(_3167_),
    .A3(_0874_),
    .ZN(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4766_ (.I(_0887_),
    .Z(_0888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4767_ (.I(_0888_),
    .Z(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4768_ (.A1(_3370_),
    .A2(_0886_),
    .B(_0889_),
    .ZN(_0890_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4769_ (.A1(_0879_),
    .A2(_0883_),
    .B(_0890_),
    .ZN(_0891_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4770_ (.I(_3355_),
    .Z(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4771_ (.I(_3176_),
    .Z(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4772_ (.I(_0875_),
    .Z(_0894_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4773_ (.A1(_0893_),
    .A2(_3285_),
    .A3(_0894_),
    .ZN(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4774_ (.I(_3176_),
    .Z(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _4775_ (.A1(_0896_),
    .A2(_3251_),
    .A3(_0894_),
    .ZN(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4776_ (.A1(_0892_),
    .A2(_0889_),
    .B(_0895_),
    .C(_0897_),
    .ZN(_0898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4777_ (.A1(_3176_),
    .A2(_0875_),
    .ZN(_0899_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4778_ (.A1(_0358_),
    .A2(_0899_),
    .ZN(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4779_ (.I(_3260_),
    .Z(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4780_ (.A1(_0901_),
    .A2(_3282_),
    .ZN(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4781_ (.A1(_0902_),
    .A2(_0899_),
    .ZN(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4782_ (.A1(_3382_),
    .A2(_0871_),
    .ZN(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _4783_ (.A1(\as2650.r0[0] ),
    .A2(_0900_),
    .B1(_0903_),
    .B2(_3342_),
    .C(_0904_),
    .ZN(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4784_ (.A1(_0891_),
    .A2(_0898_),
    .B(_0905_),
    .ZN(_0906_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4785_ (.A1(_3391_),
    .A2(_0878_),
    .B(_0906_),
    .ZN(_0907_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4786_ (.I(_0872_),
    .Z(_0908_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4787_ (.A1(_0907_),
    .A2(_0908_),
    .ZN(_0909_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4788_ (.I(_0866_),
    .Z(_0910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4789_ (.A1(_3302_),
    .A2(_0873_),
    .B(_0909_),
    .C(_0910_),
    .ZN(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4790_ (.A1(_3431_),
    .A2(_0867_),
    .B(_0911_),
    .ZN(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4791_ (.A1(_3151_),
    .A2(_3167_),
    .ZN(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4792_ (.A1(_0913_),
    .A2(_0871_),
    .ZN(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4793_ (.I(_0914_),
    .Z(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4794_ (.A1(_3151_),
    .A2(_3284_),
    .ZN(_0916_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4795_ (.A1(_0916_),
    .A2(_0871_),
    .ZN(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4796_ (.I(_0917_),
    .Z(_0918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4797_ (.A1(_3255_),
    .A2(_0663_),
    .ZN(_0919_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4798_ (.I(_0919_),
    .Z(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _4799_ (.A1(_3432_),
    .A2(_3140_),
    .A3(_3265_),
    .A4(_0920_),
    .Z(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4800_ (.A1(_3189_),
    .A2(_0894_),
    .ZN(_0922_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4801_ (.A1(_3203_),
    .A2(_0880_),
    .A3(_0654_),
    .A4(_0875_),
    .ZN(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _4802_ (.A1(_0877_),
    .A2(_0897_),
    .A3(_0922_),
    .A4(_0923_),
    .ZN(_0924_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _4803_ (.A1(_0915_),
    .A2(_0918_),
    .A3(_0921_),
    .A4(_0924_),
    .ZN(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _4804_ (.A1(_0678_),
    .A2(_0925_),
    .Z(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4805_ (.I(_0926_),
    .Z(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4806_ (.I0(_0912_),
    .I1(\as2650.r123_2[2][0] ),
    .S(_0927_),
    .Z(_0928_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4807_ (.I(_0928_),
    .Z(_0081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4808_ (.I(_0900_),
    .Z(_0929_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4809_ (.I(_0914_),
    .Z(_0930_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4810_ (.A1(_3476_),
    .A2(_0886_),
    .B(_0887_),
    .ZN(_0931_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4811_ (.A1(_3466_),
    .A2(_0882_),
    .B(_0931_),
    .ZN(_0932_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4812_ (.A1(_3461_),
    .A2(_0930_),
    .B(_0932_),
    .C(_0903_),
    .ZN(_0933_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4813_ (.A1(_3451_),
    .A2(_0903_),
    .B(_0933_),
    .ZN(_0934_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4814_ (.I(_0900_),
    .Z(_0935_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4815_ (.A1(_3482_),
    .A2(_0935_),
    .ZN(_0936_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4816_ (.I(_0876_),
    .Z(_0937_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4817_ (.A1(_0929_),
    .A2(_0934_),
    .B(_0936_),
    .C(_0937_),
    .ZN(_0938_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4818_ (.A1(_3449_),
    .A2(_0878_),
    .B(_0938_),
    .ZN(_0939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4819_ (.A1(_0908_),
    .A2(_0939_),
    .ZN(_0940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4820_ (.A1(_3492_),
    .A2(_0873_),
    .B(_0940_),
    .C(_0910_),
    .ZN(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4821_ (.A1(_3524_),
    .A2(_0867_),
    .B(_0941_),
    .ZN(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4822_ (.I0(_0942_),
    .I1(\as2650.r123_2[2][1] ),
    .S(_0927_),
    .Z(_0943_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4823_ (.I(_0943_),
    .Z(_0082_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4824_ (.I(_0866_),
    .Z(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4825_ (.A1(_3308_),
    .A2(_0894_),
    .ZN(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4826_ (.I(_0945_),
    .Z(_0946_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4827_ (.I(_0877_),
    .Z(_0947_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4828_ (.I(_0900_),
    .Z(_0948_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4829_ (.A1(_3542_),
    .A2(_0923_),
    .ZN(_0949_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4830_ (.A1(_3556_),
    .A2(_0923_),
    .B(_0914_),
    .C(_0949_),
    .ZN(_0950_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4831_ (.A1(_0346_),
    .A2(_0930_),
    .B(_0917_),
    .C(_0950_),
    .ZN(_0951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4832_ (.A1(_0892_),
    .A2(_0918_),
    .B(_0951_),
    .ZN(_0952_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4833_ (.A1(_3528_),
    .A2(_0935_),
    .ZN(_0953_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4834_ (.A1(_0948_),
    .A2(_0952_),
    .B(_0953_),
    .C(_0937_),
    .ZN(_0954_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4835_ (.A1(_3571_),
    .A2(_0947_),
    .B(_0946_),
    .C(_0954_),
    .ZN(_0955_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4836_ (.A1(_3577_),
    .A2(_0946_),
    .B(_0955_),
    .ZN(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4837_ (.A1(_0944_),
    .A2(_0956_),
    .ZN(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4838_ (.A1(_0274_),
    .A2(_0867_),
    .B(_0957_),
    .ZN(_0958_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4839_ (.I(_0926_),
    .Z(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4840_ (.I0(_0958_),
    .I1(\as2650.r123_2[2][2] ),
    .S(_0959_),
    .Z(_0960_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4841_ (.I(_0960_),
    .Z(_0083_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_2 _4842_ (.A1(_3398_),
    .A2(_0288_),
    .B1(_0311_),
    .B2(_0313_),
    .ZN(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4843_ (.I(_0917_),
    .Z(_0962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4844_ (.A1(_0345_),
    .A2(_0883_),
    .ZN(_0963_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4845_ (.A1(_0349_),
    .A2(_0883_),
    .B(_0888_),
    .C(_0963_),
    .ZN(_0964_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4846_ (.A1(_0342_),
    .A2(_0930_),
    .B(_0962_),
    .ZN(_0965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4847_ (.A1(_3546_),
    .A2(_0962_),
    .B1(_0964_),
    .B2(_0965_),
    .ZN(_0966_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4848_ (.A1(\as2650.r0[3] ),
    .A2(_0935_),
    .ZN(_0967_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4849_ (.A1(_0929_),
    .A2(_0966_),
    .B(_0967_),
    .C(_0877_),
    .ZN(_0968_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4850_ (.A1(_0331_),
    .A2(_0878_),
    .B(_0968_),
    .ZN(_0969_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4851_ (.A1(_0872_),
    .A2(_0969_),
    .ZN(_0970_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4852_ (.A1(_0325_),
    .A2(_0873_),
    .B(_0970_),
    .C(_0910_),
    .ZN(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4853_ (.A1(_0961_),
    .A2(_0867_),
    .B(_0971_),
    .ZN(_0972_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4854_ (.I0(_0972_),
    .I1(\as2650.r123_2[2][3] ),
    .S(_0959_),
    .Z(_0973_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4855_ (.I(_0973_),
    .Z(_0084_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4856_ (.I(_0393_),
    .ZN(_0974_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4857_ (.I(\as2650.r0[4] ),
    .Z(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4858_ (.I(_0346_),
    .Z(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4859_ (.A1(_3363_),
    .A2(_0874_),
    .ZN(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4860_ (.I(_0977_),
    .Z(_0978_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4861_ (.A1(_0422_),
    .A2(_0977_),
    .ZN(_0979_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4862_ (.A1(_0425_),
    .A2(_0978_),
    .B(_0888_),
    .C(_0979_),
    .ZN(_0980_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4863_ (.A1(_0463_),
    .A2(_0889_),
    .B(_0980_),
    .C(_0895_),
    .ZN(_0981_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4864_ (.A1(_0976_),
    .A2(_0895_),
    .B(_0981_),
    .C(_0897_),
    .ZN(_0982_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4865_ (.A1(_0975_),
    .A2(_0897_),
    .B(_0982_),
    .ZN(_0983_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4866_ (.A1(_0406_),
    .A2(_0937_),
    .B(_0945_),
    .ZN(_0984_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4867_ (.A1(_0947_),
    .A2(_0983_),
    .B(_0984_),
    .ZN(_0985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4868_ (.A1(_0400_),
    .A2(_0908_),
    .B(_0985_),
    .C(_0910_),
    .ZN(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _4869_ (.A1(_0974_),
    .A2(_0944_),
    .B(_0986_),
    .ZN(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4870_ (.I0(_0987_),
    .I1(\as2650.r123_2[2][4] ),
    .S(_0959_),
    .Z(_0988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4871_ (.I(_0988_),
    .Z(_0085_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4872_ (.I(_0497_),
    .Z(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4873_ (.A1(_0480_),
    .A2(_0886_),
    .B(_0888_),
    .ZN(_0990_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4874_ (.A1(_0483_),
    .A2(_0883_),
    .B(_0990_),
    .ZN(_0991_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4875_ (.A1(_0989_),
    .A2(_0915_),
    .B(_0962_),
    .C(_0991_),
    .ZN(_0992_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4876_ (.A1(_0500_),
    .A2(_0903_),
    .B(_0992_),
    .C(_0929_),
    .ZN(_0993_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4877_ (.A1(_0476_),
    .A2(_0948_),
    .B(_0993_),
    .ZN(_0994_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4878_ (.A1(_0505_),
    .A2(_0904_),
    .ZN(_0995_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4879_ (.A1(_0904_),
    .A2(_0994_),
    .B(_0995_),
    .C(_0946_),
    .ZN(_0996_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4880_ (.A1(_0475_),
    .A2(_0946_),
    .B(_0996_),
    .ZN(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4881_ (.A1(_0467_),
    .A2(_0944_),
    .ZN(_0998_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4882_ (.A1(_0944_),
    .A2(_0997_),
    .B(_0998_),
    .ZN(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4883_ (.I0(_0999_),
    .I1(\as2650.r123_2[2][5] ),
    .S(_0959_),
    .Z(_1000_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4884_ (.I(_1000_),
    .Z(_0086_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _4885_ (.A1(_0864_),
    .A2(_3272_),
    .A3(_0865_),
    .Z(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4886_ (.A1(_0556_),
    .A2(_0977_),
    .ZN(_1002_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4887_ (.A1(_0559_),
    .A2(_0978_),
    .B(_0889_),
    .C(_1002_),
    .ZN(_1003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4888_ (.A1(_3340_),
    .A2(_0930_),
    .B(_0962_),
    .ZN(_1004_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4889_ (.A1(_0463_),
    .A2(_0918_),
    .B1(_1003_),
    .B2(_1004_),
    .ZN(_1005_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4890_ (.A1(_0547_),
    .A2(_0935_),
    .ZN(_1006_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4891_ (.A1(_0929_),
    .A2(_1005_),
    .B(_1006_),
    .C(_0937_),
    .ZN(_1007_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4892_ (.A1(_0546_),
    .A2(_0878_),
    .B(_0945_),
    .C(_1007_),
    .ZN(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4893_ (.A1(_0569_),
    .A2(_0872_),
    .ZN(_1009_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4894_ (.A1(_1001_),
    .A2(_1008_),
    .A3(_1009_),
    .ZN(_1010_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4895_ (.A1(_0537_),
    .A2(_1001_),
    .B(_1010_),
    .ZN(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4896_ (.A1(\as2650.r123_2[2][6] ),
    .A2(_0927_),
    .ZN(_1012_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4897_ (.A1(_0927_),
    .A2(_1011_),
    .B(_1012_),
    .ZN(_0087_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _4898_ (.I(net8),
    .ZN(_1013_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4899_ (.I(_1013_),
    .Z(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4900_ (.A1(_1014_),
    .A2(_0978_),
    .ZN(_1015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4901_ (.A1(_0607_),
    .A2(_0978_),
    .B(_0915_),
    .C(_1015_),
    .ZN(_1016_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4902_ (.A1(_0613_),
    .A2(_0915_),
    .B(_1016_),
    .ZN(_1017_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4903_ (.A1(_0989_),
    .A2(_0918_),
    .B1(_1017_),
    .B2(_0895_),
    .ZN(_1018_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4904_ (.A1(_0617_),
    .A2(_0948_),
    .ZN(_1019_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4905_ (.A1(_0948_),
    .A2(_1018_),
    .B(_1019_),
    .C(_0947_),
    .ZN(_1020_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4906_ (.A1(_0603_),
    .A2(_0947_),
    .ZN(_1021_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4907_ (.A1(_0908_),
    .A2(_1021_),
    .ZN(_1022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _4908_ (.A1(_0623_),
    .A2(_0873_),
    .B1(_1020_),
    .B2(_1022_),
    .ZN(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4909_ (.A1(_0597_),
    .A2(_0921_),
    .ZN(_1024_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4910_ (.A1(_0921_),
    .A2(_1023_),
    .B(_1024_),
    .ZN(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _4911_ (.I0(_1025_),
    .I1(\as2650.r123_2[2][7] ),
    .S(_0926_),
    .Z(_1026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4912_ (.I(_1026_),
    .Z(_0088_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4913_ (.A1(_3170_),
    .A2(_3396_),
    .Z(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4914_ (.A1(_0675_),
    .A2(_1027_),
    .Z(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4915_ (.I(_1028_),
    .Z(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4916_ (.I(_1029_),
    .Z(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4917_ (.I(_0278_),
    .Z(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4918_ (.I(_0355_),
    .Z(_1032_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4919_ (.I(_1032_),
    .Z(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4920_ (.I(_1033_),
    .Z(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4921_ (.A1(\as2650.psl[6] ),
    .A2(_0677_),
    .Z(_1035_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _4922_ (.A1(\as2650.psl[7] ),
    .A2(_0676_),
    .Z(_1036_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4923_ (.A1(_1035_),
    .A2(_1036_),
    .ZN(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4924_ (.A1(_3137_),
    .A2(_1037_),
    .ZN(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4925_ (.A1(_1034_),
    .A2(_1038_),
    .ZN(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4926_ (.A1(_1031_),
    .A2(_1039_),
    .ZN(_1040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4927_ (.A1(_1030_),
    .A2(_1040_),
    .ZN(_1041_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4928_ (.I(_3333_),
    .Z(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4929_ (.A1(_0675_),
    .A2(_3203_),
    .ZN(_1043_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4930_ (.A1(_0310_),
    .A2(_3211_),
    .A3(_1043_),
    .ZN(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4931_ (.I(_1044_),
    .Z(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _4932_ (.A1(_1042_),
    .A2(_1045_),
    .Z(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4933_ (.A1(_3156_),
    .A2(_3178_),
    .A3(_3422_),
    .ZN(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4934_ (.A1(_3156_),
    .A2(_3547_),
    .ZN(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4935_ (.A1(_1047_),
    .A2(_1048_),
    .ZN(_1049_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4936_ (.I(_3357_),
    .Z(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4937_ (.A1(_1050_),
    .A2(_1028_),
    .ZN(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4938_ (.A1(_1049_),
    .A2(_1051_),
    .ZN(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _4939_ (.A1(_0678_),
    .A2(_1045_),
    .B(_1052_),
    .ZN(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4940_ (.A1(_3147_),
    .A2(_3219_),
    .ZN(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4941_ (.I(_1054_),
    .Z(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4942_ (.I(_1055_),
    .Z(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _4943_ (.A1(_1046_),
    .A2(_1053_),
    .B(_1056_),
    .ZN(_1057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4944_ (.A1(_1041_),
    .A2(_1057_),
    .ZN(_1058_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4945_ (.I(_0677_),
    .Z(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4946_ (.I(_1059_),
    .Z(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4947_ (.I(_1060_),
    .Z(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _4948_ (.A1(_3159_),
    .A2(_3247_),
    .ZN(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _4949_ (.A1(_0676_),
    .A2(_3158_),
    .A3(_3504_),
    .A4(_1062_),
    .ZN(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4950_ (.A1(_3209_),
    .A2(_1063_),
    .ZN(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4951_ (.I(_1064_),
    .Z(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4952_ (.I(_1065_),
    .Z(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4953_ (.I(_0893_),
    .Z(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4954_ (.A1(_3179_),
    .A2(_3173_),
    .A3(_3356_),
    .ZN(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4955_ (.I(_1068_),
    .Z(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4956_ (.A1(_3327_),
    .A2(_1069_),
    .A3(_1062_),
    .ZN(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4957_ (.I(_1070_),
    .Z(_1071_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4958_ (.A1(_1067_),
    .A2(_1071_),
    .ZN(_1072_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _4959_ (.A1(_1061_),
    .A2(_1066_),
    .B(_1072_),
    .C(_1052_),
    .ZN(_1073_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4960_ (.I(_3209_),
    .Z(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4961_ (.I(_1033_),
    .Z(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4962_ (.I(_1075_),
    .Z(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4963_ (.A1(_0868_),
    .A2(_1074_),
    .A3(_1076_),
    .A4(_1063_),
    .ZN(_1077_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4964_ (.A1(_3202_),
    .A2(_3254_),
    .ZN(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4965_ (.A1(_3218_),
    .A2(_3147_),
    .ZN(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4966_ (.A1(_1078_),
    .A2(_1079_),
    .ZN(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4967_ (.I(\as2650.halted ),
    .Z(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4968_ (.I(_3266_),
    .Z(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _4969_ (.I(_3359_),
    .Z(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4970_ (.A1(_1082_),
    .A2(_1083_),
    .ZN(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _4971_ (.A1(_0336_),
    .A2(_1068_),
    .A3(_1062_),
    .Z(_1085_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4972_ (.I(_1085_),
    .Z(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4973_ (.A1(_1081_),
    .A2(_1084_),
    .A3(_1086_),
    .ZN(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4974_ (.I(_3166_),
    .Z(_1088_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4975_ (.A1(_1088_),
    .A2(_3283_),
    .ZN(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4976_ (.I(_1089_),
    .Z(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _4977_ (.A1(_1060_),
    .A2(_1074_),
    .A3(_1063_),
    .ZN(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4978_ (.I(_1091_),
    .Z(_1092_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _4979_ (.A1(_1050_),
    .A2(_1090_),
    .A3(_1092_),
    .ZN(_1093_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4980_ (.A1(_1080_),
    .A2(_1087_),
    .A3(_1093_),
    .ZN(_1094_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _4981_ (.A1(_1058_),
    .A2(_1073_),
    .A3(_1077_),
    .A4(_1094_),
    .ZN(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _4982_ (.A1(_3206_),
    .A2(_1027_),
    .ZN(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4983_ (.I(_3236_),
    .Z(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4984_ (.A1(\as2650.r0[5] ),
    .A2(_1097_),
    .ZN(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4985_ (.I(_0481_),
    .Z(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4986_ (.I(_1099_),
    .Z(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4987_ (.I(_1100_),
    .Z(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4988_ (.I(_1101_),
    .Z(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4989_ (.I(_1102_),
    .Z(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4990_ (.I(_0357_),
    .Z(_1104_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _4991_ (.I(_1104_),
    .Z(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4992_ (.A1(_3157_),
    .A2(_3279_),
    .ZN(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _4993_ (.A1(_3174_),
    .A2(_0880_),
    .A3(_1106_),
    .ZN(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _4994_ (.I(_1107_),
    .Z(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _4995_ (.A1(_0869_),
    .A2(_1108_),
    .ZN(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4996_ (.A1(_1102_),
    .A2(_1109_),
    .ZN(_1110_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _4997_ (.A1(\as2650.psu[5] ),
    .A2(_1103_),
    .B(_1105_),
    .C(_1110_),
    .ZN(_1111_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4998_ (.A1(_1098_),
    .A2(_1111_),
    .ZN(_1112_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _4999_ (.A1(_1096_),
    .A2(_1112_),
    .ZN(_1113_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5000_ (.A1(\as2650.psu[5] ),
    .A2(_1095_),
    .ZN(_1114_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5001_ (.I(net10),
    .Z(_1115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5002_ (.I(_1115_),
    .Z(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5003_ (.A1(_1095_),
    .A2(_1113_),
    .B(_1114_),
    .C(_1116_),
    .ZN(_0089_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5004_ (.I(\as2650.psl[6] ),
    .ZN(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5005_ (.I(_1063_),
    .ZN(_1118_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5006_ (.A1(_1052_),
    .A2(_1118_),
    .A3(_1085_),
    .Z(_1119_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5007_ (.A1(_3169_),
    .A2(_3179_),
    .ZN(_1120_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5008_ (.A1(_3316_),
    .A2(_1120_),
    .ZN(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5009_ (.A1(_1070_),
    .A2(_1119_),
    .B(_1121_),
    .C(_1028_),
    .ZN(_1122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5010_ (.I(_3179_),
    .Z(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5011_ (.I(_0355_),
    .Z(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5012_ (.A1(_1123_),
    .A2(_1124_),
    .ZN(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5013_ (.I(_3362_),
    .Z(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5014_ (.I(_0663_),
    .Z(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5015_ (.A1(_1126_),
    .A2(_1127_),
    .ZN(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5016_ (.A1(_1125_),
    .A2(_1128_),
    .ZN(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5017_ (.I(_0676_),
    .Z(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5018_ (.A1(_1060_),
    .A2(_1107_),
    .ZN(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5019_ (.I(_1123_),
    .Z(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5020_ (.I(_0885_),
    .Z(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5021_ (.I(_1133_),
    .Z(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5022_ (.A1(_1132_),
    .A2(_1134_),
    .ZN(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5023_ (.A1(_1130_),
    .A2(_1131_),
    .A3(_1135_),
    .Z(_1136_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5024_ (.A1(_1122_),
    .A2(_1129_),
    .A3(_1136_),
    .ZN(_1137_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5025_ (.A1(_1132_),
    .A2(_0305_),
    .A3(_3396_),
    .ZN(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5026_ (.A1(_0305_),
    .A2(_3173_),
    .A3(_3262_),
    .A4(_3249_),
    .ZN(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5027_ (.A1(_0893_),
    .A2(_3250_),
    .A3(_1139_),
    .Z(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5028_ (.A1(_1138_),
    .A2(_1140_),
    .Z(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5029_ (.I(_0669_),
    .Z(_1142_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5030_ (.I(_1123_),
    .Z(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5031_ (.I(_1143_),
    .Z(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5032_ (.I(_3362_),
    .Z(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5033_ (.I(_1145_),
    .Z(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5034_ (.A1(_1142_),
    .A2(_1144_),
    .A3(_1031_),
    .A4(_1146_),
    .ZN(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5035_ (.A1(_0358_),
    .A2(_1141_),
    .B1(_1147_),
    .B2(_1053_),
    .ZN(_1148_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5036_ (.I(_1034_),
    .Z(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5037_ (.A1(_3254_),
    .A2(_1049_),
    .ZN(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5038_ (.A1(_3202_),
    .A2(_1096_),
    .ZN(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5039_ (.A1(_3175_),
    .A2(_3357_),
    .A3(_1150_),
    .A4(_1151_),
    .ZN(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5040_ (.I(_1146_),
    .Z(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5041_ (.I(_0355_),
    .Z(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5042_ (.A1(_3165_),
    .A2(_3262_),
    .A3(_3250_),
    .ZN(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5043_ (.A1(_3204_),
    .A2(_3212_),
    .ZN(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5044_ (.I(_3275_),
    .Z(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_2 _5045_ (.A1(_1154_),
    .A2(_1155_),
    .B1(_1156_),
    .B2(_1157_),
    .ZN(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5046_ (.A1(_1149_),
    .A2(_3285_),
    .B1(_1152_),
    .B2(_1153_),
    .C(_1158_),
    .ZN(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5047_ (.I(_0379_),
    .Z(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5048_ (.I(_3172_),
    .Z(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5049_ (.A1(_1161_),
    .A2(_1154_),
    .ZN(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5050_ (.A1(_1027_),
    .A2(_1106_),
    .ZN(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5051_ (.A1(_1161_),
    .A2(_1126_),
    .B(_1163_),
    .ZN(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5052_ (.A1(_0356_),
    .A2(_3168_),
    .ZN(_1165_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5053_ (.A1(_3207_),
    .A2(_3356_),
    .A3(_3211_),
    .ZN(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5054_ (.A1(_3204_),
    .A2(_1166_),
    .ZN(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5055_ (.A1(_0869_),
    .A2(_0358_),
    .ZN(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5056_ (.A1(_0668_),
    .A2(_0884_),
    .ZN(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5057_ (.A1(_1168_),
    .A2(_1169_),
    .B(_3152_),
    .ZN(_1170_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5058_ (.A1(_1165_),
    .A2(_1167_),
    .A3(_1170_),
    .ZN(_1171_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5059_ (.A1(_1160_),
    .A2(_1162_),
    .B(_1164_),
    .C(_1171_),
    .ZN(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5060_ (.I(_0336_),
    .Z(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5061_ (.A1(_1173_),
    .A2(_1069_),
    .A3(_1062_),
    .ZN(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5062_ (.A1(_1032_),
    .A2(_1174_),
    .ZN(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5063_ (.A1(_1081_),
    .A2(_1175_),
    .ZN(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5064_ (.A1(_0670_),
    .A2(_1079_),
    .ZN(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5065_ (.A1(_1055_),
    .A2(_1044_),
    .ZN(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5066_ (.A1(_1060_),
    .A2(_1178_),
    .ZN(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5067_ (.A1(_1173_),
    .A2(_1179_),
    .ZN(_1180_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5068_ (.A1(_1172_),
    .A2(_1176_),
    .A3(_1177_),
    .A4(_1180_),
    .Z(_1181_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5069_ (.A1(_1137_),
    .A2(_1148_),
    .A3(_1159_),
    .A4(_1181_),
    .ZN(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5070_ (.I(_3264_),
    .Z(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5071_ (.I(_0596_),
    .Z(_1184_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5072_ (.A1(_1183_),
    .A2(_1184_),
    .Z(_1185_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5073_ (.A1(_3431_),
    .A2(_3524_),
    .A3(_0274_),
    .A4(_0961_),
    .ZN(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5074_ (.A1(_0394_),
    .A2(_0467_),
    .A3(_0536_),
    .A4(_1186_),
    .ZN(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5075_ (.A1(\as2650.psl[1] ),
    .A2(_0579_),
    .ZN(_1188_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5076_ (.A1(_0514_),
    .A2(_0578_),
    .ZN(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5077_ (.A1(_3421_),
    .A2(_3401_),
    .B(_3508_),
    .ZN(_1190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5078_ (.A1(_0293_),
    .A2(_1190_),
    .B(_0288_),
    .C(_3582_),
    .ZN(_1191_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5079_ (.A1(_0375_),
    .A2(_0450_),
    .A3(_1189_),
    .ZN(_1192_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5080_ (.A1(_0296_),
    .A2(_0376_),
    .A3(_1191_),
    .B(_1192_),
    .ZN(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5081_ (.A1(_0577_),
    .A2(_0585_),
    .A3(_0586_),
    .ZN(_1194_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5082_ (.A1(_0522_),
    .A2(_1189_),
    .B(_1193_),
    .C(_1194_),
    .ZN(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5083_ (.A1(_0579_),
    .A2(_0582_),
    .B(_1188_),
    .C(_1195_),
    .ZN(_1196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5084_ (.A1(_1188_),
    .A2(_1195_),
    .B(_1196_),
    .ZN(_1197_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5085_ (.A1(_1183_),
    .A2(_1197_),
    .ZN(_1198_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5086_ (.A1(_3414_),
    .A2(_3508_),
    .A3(_0295_),
    .A4(_1192_),
    .Z(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5087_ (.A1(_0863_),
    .A2(_3236_),
    .ZN(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5088_ (.I(_1200_),
    .Z(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5089_ (.A1(_1185_),
    .A2(_1187_),
    .B1(_1198_),
    .B2(_1199_),
    .C(_1201_),
    .ZN(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5090_ (.I(_3256_),
    .Z(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5091_ (.I(_1203_),
    .Z(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5092_ (.I(_1204_),
    .Z(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5093_ (.A1(_3528_),
    .A2(_3482_),
    .A3(\as2650.r0[0] ),
    .ZN(_1206_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5094_ (.A1(\as2650.r0[6] ),
    .A2(\as2650.r0[5] ),
    .A3(\as2650.r0[4] ),
    .A4(\as2650.r0[3] ),
    .ZN(_1207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5095_ (.A1(_1206_),
    .A2(_1207_),
    .B(\as2650.r0[7] ),
    .ZN(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5096_ (.I0(_0547_),
    .I1(_1208_),
    .S(_1065_),
    .Z(_1209_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5097_ (.I(_0893_),
    .Z(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5098_ (.I(_0557_),
    .Z(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5099_ (.I(_1211_),
    .Z(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5100_ (.I(_1212_),
    .Z(_1213_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5101_ (.I(_1213_),
    .Z(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5102_ (.A1(_1173_),
    .A2(_1214_),
    .ZN(_1215_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5103_ (.A1(\as2650.psl[6] ),
    .A2(_1214_),
    .B(_1215_),
    .ZN(_1216_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5104_ (.A1(_0868_),
    .A2(_1210_),
    .A3(_1108_),
    .A4(_1216_),
    .ZN(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5105_ (.I(_1048_),
    .Z(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5106_ (.A1(_1097_),
    .A2(_1209_),
    .B(_1217_),
    .C(_1218_),
    .ZN(_1219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5107_ (.I(_3283_),
    .Z(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5108_ (.A1(_1218_),
    .A2(_0989_),
    .ZN(_1221_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5109_ (.A1(_1220_),
    .A2(_3342_),
    .A3(_0553_),
    .B(_1221_),
    .ZN(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5110_ (.I(_1088_),
    .Z(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5111_ (.A1(_1219_),
    .A2(_1222_),
    .B(_1223_),
    .ZN(_1224_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5112_ (.I(_1047_),
    .Z(_1225_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5113_ (.A1(_0500_),
    .A2(_0419_),
    .A3(_0566_),
    .ZN(_1226_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5114_ (.A1(_3529_),
    .A2(_0550_),
    .A3(_3461_),
    .A4(_0976_),
    .ZN(_1227_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5115_ (.A1(_1226_),
    .A2(_1227_),
    .B(_0613_),
    .ZN(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5116_ (.I(_3212_),
    .Z(_1229_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5117_ (.A1(_1225_),
    .A2(_1228_),
    .B(_1229_),
    .ZN(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5118_ (.I(_0611_),
    .Z(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5119_ (.I(_0884_),
    .Z(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5120_ (.A1(_1231_),
    .A2(_1232_),
    .ZN(_1233_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5121_ (.I(_0425_),
    .Z(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5122_ (.I(_0483_),
    .Z(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5123_ (.I(_0559_),
    .Z(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5124_ (.I(_0879_),
    .Z(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5125_ (.I(_3466_),
    .Z(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5126_ (.I(_3538_),
    .Z(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5127_ (.I(_1239_),
    .Z(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5128_ (.I(_1240_),
    .Z(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5129_ (.I(_0345_),
    .Z(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5130_ (.A1(_1237_),
    .A2(_1238_),
    .A3(_1241_),
    .A4(_1242_),
    .ZN(_1243_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5131_ (.A1(_1234_),
    .A2(_1235_),
    .A3(_1236_),
    .A4(_1243_),
    .ZN(_1244_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5132_ (.A1(_1224_),
    .A2(_1230_),
    .B1(_1233_),
    .B2(_1244_),
    .ZN(_1245_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5133_ (.A1(_1203_),
    .A2(_1031_),
    .A3(_3174_),
    .A4(_1074_),
    .ZN(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5134_ (.A1(_0550_),
    .A2(_1246_),
    .ZN(_1247_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5135_ (.A1(_0598_),
    .A2(_1247_),
    .ZN(_1248_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5136_ (.I(_3152_),
    .Z(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5137_ (.A1(_1143_),
    .A2(_1249_),
    .ZN(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5138_ (.A1(_1138_),
    .A2(_1208_),
    .B(_1248_),
    .C(_1250_),
    .ZN(_1251_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5139_ (.A1(_1205_),
    .A2(_1245_),
    .B(_1251_),
    .ZN(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5140_ (.A1(_1202_),
    .A2(_1252_),
    .B(_1182_),
    .ZN(_1253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5141_ (.A1(_1117_),
    .A2(_1182_),
    .B(_1253_),
    .C(_1116_),
    .ZN(_0090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5142_ (.I(\as2650.psl[7] ),
    .Z(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5143_ (.I(_1254_),
    .ZN(_1255_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5144_ (.A1(_1183_),
    .A2(_0597_),
    .B(_1198_),
    .C(_1076_),
    .ZN(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5145_ (.I(_1144_),
    .Z(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5146_ (.I(_0896_),
    .Z(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5147_ (.I(_1258_),
    .Z(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5148_ (.A1(_0617_),
    .A2(_1246_),
    .B(_1259_),
    .ZN(_1260_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5149_ (.A1(_1257_),
    .A2(_1260_),
    .ZN(_1261_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5150_ (.A1(_1247_),
    .A2(_1261_),
    .ZN(_1262_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5151_ (.I(_0884_),
    .Z(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5152_ (.I(_1263_),
    .Z(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _5153_ (.A1(_1223_),
    .A2(_0613_),
    .B(_1221_),
    .C(_1263_),
    .ZN(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5154_ (.I(_1249_),
    .Z(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5155_ (.A1(\as2650.r0[7] ),
    .A2(_1266_),
    .ZN(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5156_ (.I(_0609_),
    .Z(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5157_ (.I(net5),
    .Z(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5158_ (.I(_1269_),
    .Z(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _5159_ (.A1(_1268_),
    .A2(_3339_),
    .B1(_0342_),
    .B2(_1270_),
    .C1(_0419_),
    .C2(_1100_),
    .ZN(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5160_ (.I(_1212_),
    .Z(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5161_ (.A1(_3373_),
    .A2(_3548_),
    .B1(_3472_),
    .B2(_3464_),
    .ZN(_1273_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5162_ (.A1(_0677_),
    .A2(_0269_),
    .A3(_1068_),
    .A4(_1106_),
    .ZN(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5163_ (.A1(_3542_),
    .A2(_3546_),
    .B(_1273_),
    .C(_1274_),
    .ZN(_1275_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5164_ (.A1(_0344_),
    .A2(_0346_),
    .B1(_0566_),
    .B2(_1272_),
    .C(_1275_),
    .ZN(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5165_ (.A1(_1254_),
    .A2(_1013_),
    .B1(_3541_),
    .B2(\as2650.overflow ),
    .ZN(_1277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5166_ (.A1(_3411_),
    .A2(_3372_),
    .B1(_0344_),
    .B2(_3584_),
    .C(_1277_),
    .ZN(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5167_ (.I(\as2650.psl[1] ),
    .ZN(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5168_ (.I(_1212_),
    .Z(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5169_ (.A1(\as2650.psl[5] ),
    .A2(_0482_),
    .ZN(_1281_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5170_ (.A1(_1279_),
    .A2(_3464_),
    .B1(_1280_),
    .B2(_1117_),
    .C(_1281_),
    .ZN(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5171_ (.A1(_3253_),
    .A2(_0424_),
    .B(_1278_),
    .C(_1282_),
    .ZN(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5172_ (.I(_1043_),
    .Z(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5173_ (.A1(_0269_),
    .A2(_1069_),
    .ZN(_1285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5174_ (.A1(_1059_),
    .A2(_1283_),
    .B(_1284_),
    .C(_1285_),
    .ZN(_1286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5175_ (.A1(_1271_),
    .A2(_1276_),
    .B(_1286_),
    .ZN(_1287_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5176_ (.I(\as2650.psu[4] ),
    .ZN(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5177_ (.I(_1270_),
    .Z(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5178_ (.I(net24),
    .ZN(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5179_ (.I(_3373_),
    .ZN(_1291_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5180_ (.I(_3464_),
    .ZN(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5181_ (.A1(\as2650.psu[0] ),
    .A2(_1291_),
    .B1(_1292_),
    .B2(\as2650.psu[1] ),
    .ZN(_1293_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5182_ (.A1(_1288_),
    .A2(_1289_),
    .B1(_1214_),
    .B2(_1290_),
    .C(_1293_),
    .ZN(_1294_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5183_ (.I(\as2650.psu[7] ),
    .ZN(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5184_ (.I(\as2650.psu[5] ),
    .ZN(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5185_ (.I(net4),
    .ZN(_1297_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5186_ (.I(_1297_),
    .Z(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5187_ (.A1(\as2650.psu[2] ),
    .A2(_3542_),
    .B1(_1298_),
    .B2(\as2650.psu[3] ),
    .ZN(_1299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5188_ (.A1(_1295_),
    .A2(_1268_),
    .B1(_1101_),
    .B2(_1296_),
    .C(_1299_),
    .ZN(_1300_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5189_ (.A1(_1059_),
    .A2(_1284_),
    .ZN(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5190_ (.A1(_1161_),
    .A2(_3506_),
    .A3(_1301_),
    .ZN(_1302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5191_ (.A1(_1294_),
    .A2(_1300_),
    .B(_1302_),
    .ZN(_1303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5192_ (.A1(_3138_),
    .A2(_1045_),
    .B(_1287_),
    .C(_1303_),
    .ZN(_1304_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5193_ (.A1(_1254_),
    .A2(_0611_),
    .A3(_0678_),
    .A4(_1108_),
    .ZN(_1305_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5194_ (.A1(_1046_),
    .A2(_1304_),
    .A3(_1305_),
    .ZN(_1306_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5195_ (.I(_0611_),
    .Z(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5196_ (.A1(_1042_),
    .A2(_1045_),
    .ZN(_1308_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5197_ (.A1(_1255_),
    .A2(_1307_),
    .A3(_1308_),
    .ZN(_1309_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5198_ (.I(_1033_),
    .Z(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5199_ (.A1(_1306_),
    .A2(_1309_),
    .B(_1310_),
    .ZN(_1311_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5200_ (.I(_1089_),
    .Z(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5201_ (.A1(_1267_),
    .A2(_1311_),
    .B(_1312_),
    .ZN(_1313_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5202_ (.A1(_1231_),
    .A2(_1264_),
    .B1(_1265_),
    .B2(_1313_),
    .ZN(_1314_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5203_ (.A1(_1256_),
    .A2(_1262_),
    .B1(_1314_),
    .B2(_1205_),
    .ZN(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5204_ (.A1(_1182_),
    .A2(_1315_),
    .ZN(_1316_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5205_ (.A1(_1255_),
    .A2(_1182_),
    .B(_1316_),
    .C(_1116_),
    .ZN(_0091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5206_ (.I(_3147_),
    .Z(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5207_ (.A1(_1317_),
    .A2(_3304_),
    .ZN(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5208_ (.I(_1318_),
    .Z(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5209_ (.A1(_1237_),
    .A2(_1319_),
    .ZN(_1320_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5210_ (.I(_3274_),
    .Z(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5211_ (.I(_1317_),
    .Z(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5212_ (.A1(_0610_),
    .A2(_1126_),
    .ZN(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5213_ (.I(_0675_),
    .Z(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5214_ (.A1(_1324_),
    .A2(_0672_),
    .ZN(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5215_ (.I(_1325_),
    .Z(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5216_ (.I(_1326_),
    .Z(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5217_ (.A1(_0683_),
    .A2(_1327_),
    .B(_0653_),
    .ZN(_1328_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5218_ (.A1(_1321_),
    .A2(_1322_),
    .A3(_1323_),
    .A4(_1328_),
    .ZN(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5219_ (.A1(_1329_),
    .A2(_1319_),
    .Z(_1330_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5220_ (.I(_1329_),
    .Z(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5221_ (.A1(_1061_),
    .A2(_1331_),
    .ZN(_1332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5222_ (.A1(_1320_),
    .A2(_1330_),
    .B(_1332_),
    .ZN(_0092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5223_ (.I(_1238_),
    .Z(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5224_ (.A1(_1333_),
    .A2(_1319_),
    .ZN(_1334_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5225_ (.A1(_1130_),
    .A2(_1329_),
    .ZN(_1335_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5226_ (.A1(_1330_),
    .A2(_1334_),
    .B(_1335_),
    .ZN(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5227_ (.I(_3157_),
    .Z(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5228_ (.I(_1336_),
    .Z(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5229_ (.I(_1337_),
    .Z(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5230_ (.A1(_1082_),
    .A2(_1321_),
    .A3(_1322_),
    .A4(_3434_),
    .ZN(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5231_ (.A1(_1241_),
    .A2(_1339_),
    .ZN(_1340_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5232_ (.A1(_1338_),
    .A2(_1331_),
    .B(_1340_),
    .ZN(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5233_ (.A1(_1336_),
    .A2(_0680_),
    .ZN(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5234_ (.I(_1341_),
    .Z(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5235_ (.I(_1342_),
    .Z(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5236_ (.I(_1343_),
    .Z(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5237_ (.I(_1344_),
    .Z(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5238_ (.A1(_1345_),
    .A2(_1329_),
    .B(_1031_),
    .ZN(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5239_ (.A1(_1103_),
    .A2(_1339_),
    .ZN(_1347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5240_ (.A1(_1330_),
    .A2(_1346_),
    .B(_1347_),
    .ZN(_0095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5241_ (.I(_1214_),
    .Z(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5242_ (.I(_1348_),
    .Z(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5243_ (.A1(_1349_),
    .A2(_1339_),
    .ZN(_1350_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5244_ (.A1(_3504_),
    .A2(_1331_),
    .B(_1350_),
    .ZN(_0096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5245_ (.I(_1307_),
    .Z(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5246_ (.A1(_1351_),
    .A2(_1339_),
    .ZN(_1352_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5247_ (.A1(_3356_),
    .A2(_1331_),
    .B(_1352_),
    .ZN(_0097_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5248_ (.A1(_0689_),
    .A2(_0782_),
    .ZN(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5249_ (.I(_1353_),
    .Z(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5250_ (.I(_1354_),
    .Z(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5251_ (.I(_1353_),
    .Z(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5252_ (.A1(\as2650.stack[6][0] ),
    .A2(_1356_),
    .ZN(_1357_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5253_ (.A1(_0835_),
    .A2(_1355_),
    .B(_1357_),
    .ZN(_0098_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5254_ (.A1(\as2650.stack[6][1] ),
    .A2(_1356_),
    .ZN(_1358_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5255_ (.A1(_0841_),
    .A2(_1355_),
    .B(_1358_),
    .ZN(_0099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5256_ (.A1(\as2650.stack[6][2] ),
    .A2(_1356_),
    .ZN(_1359_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5257_ (.A1(_0813_),
    .A2(_1355_),
    .B(_1359_),
    .ZN(_0100_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5258_ (.A1(\as2650.stack[6][3] ),
    .A2(_1356_),
    .ZN(_1360_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5259_ (.A1(_0815_),
    .A2(_1355_),
    .B(_1360_),
    .ZN(_0101_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5260_ (.I(_1354_),
    .Z(_1361_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5261_ (.I(_1353_),
    .Z(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5262_ (.A1(\as2650.stack[6][4] ),
    .A2(_1362_),
    .ZN(_1363_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5263_ (.A1(_0817_),
    .A2(_1361_),
    .B(_1363_),
    .ZN(_0102_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5264_ (.A1(\as2650.stack[6][5] ),
    .A2(_1362_),
    .ZN(_1364_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5265_ (.A1(_0821_),
    .A2(_1361_),
    .B(_1364_),
    .ZN(_0103_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5266_ (.A1(\as2650.stack[6][6] ),
    .A2(_1362_),
    .ZN(_1365_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5267_ (.A1(_0823_),
    .A2(_1361_),
    .B(_1365_),
    .ZN(_0104_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5268_ (.A1(\as2650.stack[6][7] ),
    .A2(_1362_),
    .ZN(_1366_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5269_ (.A1(_0850_),
    .A2(_1361_),
    .B(_1366_),
    .ZN(_0105_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5270_ (.I0(_0852_),
    .I1(\as2650.stack[6][8] ),
    .S(_1354_),
    .Z(_1367_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5271_ (.I(_1367_),
    .Z(_0106_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5272_ (.I(_1354_),
    .Z(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5273_ (.I(_1353_),
    .Z(_1369_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5274_ (.A1(\as2650.stack[6][9] ),
    .A2(_1369_),
    .ZN(_1370_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5275_ (.A1(_0827_),
    .A2(_1368_),
    .B(_1370_),
    .ZN(_0107_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5276_ (.A1(\as2650.stack[6][10] ),
    .A2(_1369_),
    .ZN(_1371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5277_ (.A1(_0831_),
    .A2(_1368_),
    .B(_1371_),
    .ZN(_0108_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5278_ (.A1(\as2650.stack[6][11] ),
    .A2(_1369_),
    .ZN(_1372_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5279_ (.A1(_0858_),
    .A2(_1368_),
    .B(_1372_),
    .ZN(_0109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5280_ (.A1(\as2650.stack[6][12] ),
    .A2(_1369_),
    .ZN(_1373_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5281_ (.A1(_0860_),
    .A2(_1368_),
    .B(_1373_),
    .ZN(_0110_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5282_ (.A1(_1061_),
    .A2(_0925_),
    .ZN(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5283_ (.I(_1374_),
    .Z(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5284_ (.I0(\as2650.r123_2[1][0] ),
    .I1(_0912_),
    .S(_1375_),
    .Z(_1376_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5285_ (.I(_1376_),
    .Z(_0111_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5286_ (.I0(\as2650.r123_2[1][1] ),
    .I1(_0942_),
    .S(_1375_),
    .Z(_1377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5287_ (.I(_1377_),
    .Z(_0112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5288_ (.I(_1374_),
    .Z(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5289_ (.I0(\as2650.r123_2[1][2] ),
    .I1(_0958_),
    .S(_1378_),
    .Z(_1379_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5290_ (.I(_1379_),
    .Z(_0113_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5291_ (.I0(\as2650.r123_2[1][3] ),
    .I1(_0972_),
    .S(_1378_),
    .Z(_1380_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5292_ (.I(_1380_),
    .Z(_0114_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5293_ (.I0(\as2650.r123_2[1][4] ),
    .I1(_0987_),
    .S(_1378_),
    .Z(_1381_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5294_ (.I(_1381_),
    .Z(_0115_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5295_ (.I(_1378_),
    .Z(_1382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5296_ (.A1(_0999_),
    .A2(_1382_),
    .ZN(_1383_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5297_ (.A1(_0413_),
    .A2(_1382_),
    .B(_1383_),
    .ZN(_0116_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5298_ (.I(_1011_),
    .ZN(_1384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5299_ (.A1(_1384_),
    .A2(_1375_),
    .ZN(_1385_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5300_ (.A1(_0492_),
    .A2(_1382_),
    .B(_1385_),
    .ZN(_0117_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5301_ (.A1(_1025_),
    .A2(_1375_),
    .ZN(_1386_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5302_ (.A1(_3328_),
    .A2(_1382_),
    .B(_1386_),
    .ZN(_0118_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5303_ (.I(\as2650.r123[3][0] ),
    .Z(_1387_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5304_ (.I(_1387_),
    .Z(_0119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5305_ (.I(\as2650.r123[3][1] ),
    .Z(_1388_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5306_ (.I(_1388_),
    .Z(_0120_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5307_ (.I(\as2650.r123[3][2] ),
    .Z(_1389_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5308_ (.I(_1389_),
    .Z(_0121_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5309_ (.I(\as2650.r123[3][3] ),
    .Z(_1390_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5310_ (.I(_1390_),
    .Z(_0122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5311_ (.I(\as2650.r123[3][4] ),
    .Z(_1391_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5312_ (.I(_1391_),
    .Z(_0123_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5313_ (.I(\as2650.r123[3][5] ),
    .Z(_1392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5314_ (.I(_1392_),
    .Z(_0124_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5315_ (.I(\as2650.r123[3][6] ),
    .Z(_1393_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5316_ (.I(_1393_),
    .Z(_0125_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5317_ (.I(\as2650.r123[3][7] ),
    .Z(_1394_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5318_ (.I(_1394_),
    .Z(_0126_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5319_ (.A1(_0689_),
    .A2(_0806_),
    .ZN(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5320_ (.I(_1395_),
    .Z(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5321_ (.I(_1396_),
    .Z(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5322_ (.I(_1395_),
    .Z(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5323_ (.A1(\as2650.stack[5][0] ),
    .A2(_1398_),
    .ZN(_1399_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5324_ (.A1(_0835_),
    .A2(_1397_),
    .B(_1399_),
    .ZN(_0127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5325_ (.A1(\as2650.stack[5][1] ),
    .A2(_1398_),
    .ZN(_1400_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5326_ (.A1(_0841_),
    .A2(_1397_),
    .B(_1400_),
    .ZN(_0128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5327_ (.A1(\as2650.stack[5][2] ),
    .A2(_1398_),
    .ZN(_1401_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5328_ (.A1(_0813_),
    .A2(_1397_),
    .B(_1401_),
    .ZN(_0129_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5329_ (.A1(\as2650.stack[5][3] ),
    .A2(_1398_),
    .ZN(_1402_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5330_ (.A1(_0815_),
    .A2(_1397_),
    .B(_1402_),
    .ZN(_0130_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5331_ (.I(_1396_),
    .Z(_1403_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5332_ (.I(_1395_),
    .Z(_1404_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5333_ (.A1(\as2650.stack[5][4] ),
    .A2(_1404_),
    .ZN(_1405_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5334_ (.A1(_0817_),
    .A2(_1403_),
    .B(_1405_),
    .ZN(_0131_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5335_ (.A1(\as2650.stack[5][5] ),
    .A2(_1404_),
    .ZN(_1406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5336_ (.A1(_0821_),
    .A2(_1403_),
    .B(_1406_),
    .ZN(_0132_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5337_ (.A1(\as2650.stack[5][6] ),
    .A2(_1404_),
    .ZN(_1407_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5338_ (.A1(_0823_),
    .A2(_1403_),
    .B(_1407_),
    .ZN(_0133_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5339_ (.A1(\as2650.stack[5][7] ),
    .A2(_1404_),
    .ZN(_1408_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5340_ (.A1(_0850_),
    .A2(_1403_),
    .B(_1408_),
    .ZN(_0134_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5341_ (.I0(_0852_),
    .I1(\as2650.stack[5][8] ),
    .S(_1396_),
    .Z(_1409_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5342_ (.I(_1409_),
    .Z(_0135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5343_ (.I(_1396_),
    .Z(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5344_ (.I(_1395_),
    .Z(_1411_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5345_ (.A1(\as2650.stack[5][9] ),
    .A2(_1411_),
    .ZN(_1412_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5346_ (.A1(_0827_),
    .A2(_1410_),
    .B(_1412_),
    .ZN(_0136_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5347_ (.A1(\as2650.stack[5][10] ),
    .A2(_1411_),
    .ZN(_1413_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5348_ (.A1(_0831_),
    .A2(_1410_),
    .B(_1413_),
    .ZN(_0137_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5349_ (.A1(\as2650.stack[5][11] ),
    .A2(_1411_),
    .ZN(_1414_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5350_ (.A1(_0858_),
    .A2(_1410_),
    .B(_1414_),
    .ZN(_0138_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5351_ (.A1(\as2650.stack[5][12] ),
    .A2(_1411_),
    .ZN(_1415_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5352_ (.A1(_0860_),
    .A2(_1410_),
    .B(_1415_),
    .ZN(_0139_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5353_ (.I(_3270_),
    .Z(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5354_ (.I(_1416_),
    .Z(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5355_ (.I(_1417_),
    .Z(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5356_ (.A1(_3266_),
    .A2(_0656_),
    .ZN(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5357_ (.I(_1419_),
    .Z(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5358_ (.A1(_1336_),
    .A2(_0671_),
    .ZN(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5359_ (.I(_1421_),
    .Z(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5360_ (.I(_1422_),
    .Z(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5361_ (.I(_1423_),
    .Z(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5362_ (.A1(_1418_),
    .A2(_1420_),
    .A3(_1424_),
    .ZN(_1425_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5363_ (.I(_1157_),
    .Z(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5364_ (.A1(_0669_),
    .A2(_1343_),
    .ZN(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5365_ (.A1(_1426_),
    .A2(_1427_),
    .ZN(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5366_ (.I(_1416_),
    .Z(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5367_ (.I(_0681_),
    .Z(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5368_ (.I(_1430_),
    .Z(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5369_ (.A1(_3169_),
    .A2(_3151_),
    .A3(_0672_),
    .ZN(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5370_ (.I(_1324_),
    .Z(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5371_ (.I(_0668_),
    .Z(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5372_ (.I(_1054_),
    .Z(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5373_ (.I(_0672_),
    .Z(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5374_ (.A1(_1433_),
    .A2(_1434_),
    .A3(_1435_),
    .A4(_1436_),
    .ZN(_1437_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5375_ (.A1(_1429_),
    .A2(_1431_),
    .B(_1432_),
    .C(_1437_),
    .ZN(_1438_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5376_ (.I(_0668_),
    .Z(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5377_ (.A1(_1027_),
    .A2(_1038_),
    .Z(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5378_ (.A1(_1124_),
    .A2(_1284_),
    .ZN(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5379_ (.A1(_1440_),
    .A2(_1441_),
    .ZN(_1442_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5380_ (.A1(_1151_),
    .A2(_1342_),
    .ZN(_1443_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5381_ (.I(_1081_),
    .Z(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5382_ (.A1(_1434_),
    .A2(_0667_),
    .B(_1443_),
    .C(_1444_),
    .ZN(_1445_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5383_ (.A1(_1439_),
    .A2(_1266_),
    .B(_1442_),
    .C(_1445_),
    .ZN(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5384_ (.A1(_1438_),
    .A2(_1446_),
    .Z(_1447_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5385_ (.A1(_3266_),
    .A2(_0656_),
    .Z(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5386_ (.A1(_0660_),
    .A2(_1448_),
    .ZN(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5387_ (.A1(_0356_),
    .A2(_1133_),
    .A3(_0673_),
    .A4(_1449_),
    .ZN(_1450_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5388_ (.I(_3181_),
    .Z(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5389_ (.A1(_1451_),
    .A2(_0662_),
    .ZN(_1452_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5390_ (.I(_1452_),
    .Z(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5391_ (.A1(_0658_),
    .A2(_1453_),
    .A3(_0673_),
    .ZN(_1454_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5392_ (.I(_3204_),
    .Z(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5393_ (.A1(_1450_),
    .A2(_1454_),
    .B(_1455_),
    .ZN(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5394_ (.A1(_1425_),
    .A2(_1428_),
    .B(_1447_),
    .C(_1456_),
    .ZN(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5395_ (.I(_1457_),
    .Z(_1458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5396_ (.I(_3238_),
    .Z(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5397_ (.I(_1459_),
    .Z(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5398_ (.I(_1460_),
    .Z(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5399_ (.A1(_0751_),
    .A2(_1458_),
    .B(_1461_),
    .ZN(_1462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5400_ (.A1(_0751_),
    .A2(_1458_),
    .B(_1462_),
    .ZN(_0140_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5401_ (.I(_1142_),
    .Z(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5402_ (.A1(_0651_),
    .A2(_0755_),
    .B(_1463_),
    .ZN(_1464_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5403_ (.I(_1439_),
    .Z(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5404_ (.I(_1465_),
    .Z(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5405_ (.A1(_1466_),
    .A2(_0651_),
    .A3(_0755_),
    .Z(_1467_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5406_ (.A1(_1464_),
    .A2(_1467_),
    .ZN(_1468_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5407_ (.I(_1459_),
    .Z(_1469_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5408_ (.I(_1469_),
    .Z(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5409_ (.A1(\as2650.stack_ptr[1] ),
    .A2(_1457_),
    .B(_1470_),
    .ZN(_1471_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5410_ (.A1(_1458_),
    .A2(_1468_),
    .B(_1471_),
    .ZN(_0141_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5411_ (.A1(\as2650.stack_ptr[2] ),
    .A2(_0648_),
    .Z(_1472_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5412_ (.I(_1472_),
    .Z(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5413_ (.A1(_1464_),
    .A2(_1473_),
    .Z(_1474_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5414_ (.A1(_0652_),
    .A2(_1457_),
    .B(_1470_),
    .ZN(_1475_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5415_ (.A1(_1458_),
    .A2(_1474_),
    .B(_1475_),
    .ZN(_0142_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5416_ (.A1(_1130_),
    .A2(_0925_),
    .ZN(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5417_ (.I(_1476_),
    .Z(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5418_ (.I0(\as2650.r123_2[0][0] ),
    .I1(_0912_),
    .S(_1477_),
    .Z(_1478_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5419_ (.I(_1478_),
    .Z(_0143_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5420_ (.I0(\as2650.r123_2[0][1] ),
    .I1(_0942_),
    .S(_1477_),
    .Z(_1479_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5421_ (.I(_1479_),
    .Z(_0144_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5422_ (.I(_1476_),
    .Z(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5423_ (.I0(\as2650.r123_2[0][2] ),
    .I1(_0958_),
    .S(_1480_),
    .Z(_1481_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5424_ (.I(_1481_),
    .Z(_0145_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5425_ (.I0(\as2650.r123_2[0][3] ),
    .I1(_0972_),
    .S(_1480_),
    .Z(_1482_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5426_ (.I(_1482_),
    .Z(_0146_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5427_ (.I0(\as2650.r123_2[0][4] ),
    .I1(_0987_),
    .S(_1480_),
    .Z(_1483_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5428_ (.I(_1483_),
    .Z(_0147_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5429_ (.I(_1480_),
    .Z(_1484_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5430_ (.A1(_0999_),
    .A2(_1484_),
    .ZN(_1485_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5431_ (.A1(_0410_),
    .A2(_1484_),
    .B(_1485_),
    .ZN(_0148_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5432_ (.A1(_1384_),
    .A2(_1477_),
    .ZN(_1486_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5433_ (.A1(_0489_),
    .A2(_1484_),
    .B(_1486_),
    .ZN(_0149_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5434_ (.A1(_1025_),
    .A2(_1477_),
    .ZN(_1487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5435_ (.A1(_3334_),
    .A2(_1484_),
    .B(_1487_),
    .ZN(_0150_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5436_ (.I(_1291_),
    .Z(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5437_ (.I(_0660_),
    .Z(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5438_ (.A1(_1489_),
    .A2(_1419_),
    .ZN(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5439_ (.A1(_1127_),
    .A2(_1490_),
    .ZN(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5440_ (.A1(_0661_),
    .A2(_0684_),
    .ZN(_1492_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5441_ (.A1(_0660_),
    .A2(_1492_),
    .ZN(_1493_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5442_ (.A1(_1054_),
    .A2(_1493_),
    .ZN(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5443_ (.I(_3142_),
    .Z(_1495_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5444_ (.A1(_3215_),
    .A2(_3216_),
    .A3(_3218_),
    .A4(\as2650.cycle[0] ),
    .ZN(_1496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5445_ (.I(_1496_),
    .Z(_1497_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5446_ (.A1(_3224_),
    .A2(_1495_),
    .A3(_1497_),
    .Z(_1498_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5447_ (.A1(_1419_),
    .A2(_1498_),
    .ZN(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5448_ (.A1(_3182_),
    .A2(_3183_),
    .A3(_3225_),
    .ZN(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5449_ (.A1(\as2650.cycle[6] ),
    .A2(_1495_),
    .A3(_1496_),
    .ZN(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5450_ (.A1(_3224_),
    .A2(_1501_),
    .ZN(_1502_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5451_ (.A1(_1500_),
    .A2(_1502_),
    .ZN(_1503_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5452_ (.A1(_1494_),
    .A2(_1499_),
    .A3(_1503_),
    .Z(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5453_ (.A1(_1491_),
    .A2(_1504_),
    .B(_1200_),
    .ZN(_1505_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5454_ (.I(_0670_),
    .Z(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5455_ (.A1(_3271_),
    .A2(_1449_),
    .ZN(_1507_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5456_ (.A1(_1133_),
    .A2(_1506_),
    .A3(_1430_),
    .A4(_1507_),
    .ZN(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5457_ (.A1(_3221_),
    .A2(_0681_),
    .ZN(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5458_ (.A1(_1492_),
    .A2(_1509_),
    .ZN(_1510_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5459_ (.I(_1342_),
    .Z(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5460_ (.I(_1493_),
    .Z(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5461_ (.I(_1512_),
    .Z(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5462_ (.I(_1506_),
    .Z(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5463_ (.A1(_1513_),
    .A2(_1514_),
    .A3(_1343_),
    .ZN(_1515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5464_ (.I(_1120_),
    .Z(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5465_ (.I(_1079_),
    .Z(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5466_ (.I(_1517_),
    .Z(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5467_ (.I(_3226_),
    .Z(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5468_ (.A1(_3172_),
    .A2(_1519_),
    .ZN(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5469_ (.A1(_3434_),
    .A2(_1516_),
    .A3(_1518_),
    .A4(_1520_),
    .ZN(_1521_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5470_ (.A1(_1075_),
    .A2(_1511_),
    .A3(_1515_),
    .A4(_1521_),
    .ZN(_1522_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5471_ (.I(_3362_),
    .Z(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5472_ (.I(_0679_),
    .Z(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5473_ (.I(_0680_),
    .Z(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5474_ (.A1(_3207_),
    .A2(_1523_),
    .A3(_1524_),
    .A4(_1525_),
    .ZN(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5475_ (.I(\as2650.cycle[6] ),
    .Z(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5476_ (.I(_1527_),
    .ZN(_1528_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5477_ (.A1(_1528_),
    .A2(_1498_),
    .ZN(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5478_ (.I(_1529_),
    .Z(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5479_ (.A1(_0864_),
    .A2(_1530_),
    .ZN(_1531_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5480_ (.I(_1449_),
    .ZN(_1532_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _5481_ (.A1(_1523_),
    .A2(_1532_),
    .B(_3255_),
    .ZN(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5482_ (.A1(_1522_),
    .A2(_1526_),
    .A3(_1531_),
    .A4(_1533_),
    .ZN(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5483_ (.A1(_1505_),
    .A2(_1508_),
    .A3(_1510_),
    .A4(_1534_),
    .ZN(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5484_ (.I(_1535_),
    .Z(_1536_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5485_ (.I(\as2650.addr_buff[0] ),
    .Z(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5486_ (.I(_1535_),
    .Z(_1538_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5487_ (.A1(_1537_),
    .A2(_1538_),
    .ZN(_1539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5488_ (.A1(_1488_),
    .A2(_1536_),
    .B(_1539_),
    .ZN(_0151_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5489_ (.I(\as2650.addr_buff[1] ),
    .Z(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5490_ (.A1(_1540_),
    .A2(_1538_),
    .ZN(_1541_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5491_ (.A1(_1292_),
    .A2(_1536_),
    .B(_1541_),
    .ZN(_0152_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5492_ (.I(\as2650.addr_buff[2] ),
    .Z(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5493_ (.A1(_1542_),
    .A2(_1538_),
    .ZN(_1543_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5494_ (.A1(_3543_),
    .A2(_1536_),
    .B(_1543_),
    .ZN(_0153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5495_ (.I(_1298_),
    .Z(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5496_ (.I(\as2650.addr_buff[3] ),
    .Z(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5497_ (.A1(_1545_),
    .A2(_1538_),
    .ZN(_1546_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5498_ (.A1(_1544_),
    .A2(_1536_),
    .B(_1546_),
    .ZN(_0154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5499_ (.I(_1535_),
    .Z(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5500_ (.I(\as2650.addr_buff[4] ),
    .Z(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5501_ (.I(_1535_),
    .Z(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5502_ (.A1(_1548_),
    .A2(_1549_),
    .ZN(_1550_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5503_ (.A1(_1234_),
    .A2(_1547_),
    .B(_1550_),
    .ZN(_0155_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5504_ (.A1(_3228_),
    .A2(_1549_),
    .ZN(_1551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5505_ (.A1(_1235_),
    .A2(_1547_),
    .B(_1551_),
    .ZN(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5506_ (.A1(_3229_),
    .A2(_1549_),
    .ZN(_1552_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5507_ (.A1(_1236_),
    .A2(_1547_),
    .B(_1552_),
    .ZN(_0157_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5508_ (.I(_1014_),
    .Z(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5509_ (.I(_1553_),
    .Z(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5510_ (.I(_0659_),
    .Z(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5511_ (.A1(_1555_),
    .A2(_1549_),
    .ZN(_1556_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5512_ (.A1(_1554_),
    .A2(_1547_),
    .B(_1556_),
    .ZN(_0158_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5513_ (.A1(_0661_),
    .A2(_3359_),
    .ZN(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5514_ (.I(_1557_),
    .Z(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5515_ (.A1(_1051_),
    .A2(_1120_),
    .ZN(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5516_ (.A1(_1524_),
    .A2(_1558_),
    .A3(_1156_),
    .A4(_1559_),
    .ZN(_1560_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5517_ (.A1(_0920_),
    .A2(_1162_),
    .A3(_1560_),
    .Z(_1561_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5518_ (.I(_3271_),
    .Z(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5519_ (.A1(_1074_),
    .A2(_1050_),
    .ZN(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _5520_ (.A1(_1083_),
    .A2(_1562_),
    .A3(_1563_),
    .ZN(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5521_ (.A1(_1448_),
    .A2(_1129_),
    .ZN(_1565_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5522_ (.I(_0896_),
    .Z(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5523_ (.I(_1566_),
    .Z(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5524_ (.I(_1444_),
    .Z(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5525_ (.A1(_1567_),
    .A2(_1166_),
    .B(_1164_),
    .C(_1568_),
    .ZN(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5526_ (.A1(_1565_),
    .A2(_1569_),
    .ZN(_1570_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5527_ (.A1(_1561_),
    .A2(_1564_),
    .A3(_1570_),
    .ZN(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5528_ (.I(_1257_),
    .Z(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5529_ (.A1(_1572_),
    .A2(_1449_),
    .B(_1135_),
    .ZN(_1573_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5530_ (.A1(net21),
    .A2(_1571_),
    .ZN(_1574_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5531_ (.I(_3438_),
    .Z(_1575_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5532_ (.I(_1575_),
    .Z(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5533_ (.A1(_1571_),
    .A2(_1573_),
    .B(_1574_),
    .C(_1576_),
    .ZN(_0159_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5534_ (.I(_1444_),
    .Z(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5535_ (.I(_1076_),
    .Z(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5536_ (.A1(_3203_),
    .A2(_1050_),
    .ZN(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5537_ (.A1(_1577_),
    .A2(_1578_),
    .A3(_1579_),
    .ZN(_1580_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5538_ (.A1(net45),
    .A2(_1580_),
    .B(_1470_),
    .ZN(_1581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5539_ (.A1(_3504_),
    .A2(_1580_),
    .B(_1581_),
    .ZN(_0160_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5540_ (.I(net20),
    .ZN(_1582_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5541_ (.I(_1516_),
    .Z(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5542_ (.A1(_1145_),
    .A2(_1167_),
    .B1(_1163_),
    .B2(_1518_),
    .ZN(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5543_ (.A1(_1051_),
    .A2(_1080_),
    .ZN(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5544_ (.A1(_1577_),
    .A2(_1318_),
    .ZN(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5545_ (.I(_1455_),
    .Z(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5546_ (.A1(_1451_),
    .A2(_1557_),
    .ZN(_1588_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5547_ (.I(_1588_),
    .Z(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5548_ (.A1(_1587_),
    .A2(_1589_),
    .ZN(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5549_ (.A1(_1203_),
    .A2(_1518_),
    .ZN(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5550_ (.A1(_1322_),
    .A2(_1169_),
    .B(_1590_),
    .C(_1591_),
    .ZN(_1592_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5551_ (.A1(_1585_),
    .A2(_1586_),
    .A3(_1592_),
    .ZN(_1593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5552_ (.A1(_1583_),
    .A2(_1564_),
    .B(_1584_),
    .C(_1593_),
    .ZN(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5553_ (.I(_1115_),
    .Z(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5554_ (.A1(_3149_),
    .A2(_1594_),
    .B(_1595_),
    .ZN(_1596_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5555_ (.A1(_1582_),
    .A2(_1594_),
    .B(_1596_),
    .ZN(_0161_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5556_ (.A1(_3305_),
    .A2(_1504_),
    .ZN(_1597_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5557_ (.A1(_0683_),
    .A2(_3274_),
    .A3(_0685_),
    .ZN(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5558_ (.A1(_0862_),
    .A2(_1083_),
    .ZN(_1599_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5559_ (.A1(_1598_),
    .A2(_1499_),
    .A3(_1599_),
    .ZN(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5560_ (.A1(_1597_),
    .A2(_1600_),
    .ZN(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5561_ (.A1(_1140_),
    .A2(_1601_),
    .ZN(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5562_ (.A1(_1069_),
    .A2(_1037_),
    .B(_1440_),
    .ZN(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5563_ (.A1(_1432_),
    .A2(_1603_),
    .ZN(_1604_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5564_ (.A1(_1175_),
    .A2(_1604_),
    .ZN(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5565_ (.A1(_1047_),
    .A2(_1080_),
    .B(_1081_),
    .ZN(_1606_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5566_ (.A1(_1083_),
    .A2(_1524_),
    .A3(_1341_),
    .B(_1606_),
    .ZN(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _5567_ (.A1(_1258_),
    .A2(_1066_),
    .B1(_1516_),
    .B2(_1564_),
    .C(_1607_),
    .ZN(_1608_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5568_ (.A1(_1048_),
    .A2(_1177_),
    .ZN(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5569_ (.A1(_1558_),
    .A2(_1152_),
    .ZN(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5570_ (.A1(_1608_),
    .A2(_1609_),
    .A3(_1610_),
    .ZN(_1611_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5571_ (.A1(_3214_),
    .A2(_1497_),
    .ZN(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5572_ (.I(_1612_),
    .Z(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5573_ (.A1(_1075_),
    .A2(_1514_),
    .A3(_1436_),
    .A4(_1613_),
    .ZN(_1614_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5574_ (.A1(_1323_),
    .A2(_1325_),
    .B(_1533_),
    .ZN(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5575_ (.A1(_1144_),
    .A2(_1429_),
    .B1(_1520_),
    .B2(_1555_),
    .C(_1318_),
    .ZN(_1616_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5576_ (.A1(_1527_),
    .A2(_1495_),
    .A3(_1497_),
    .Z(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5577_ (.A1(_1161_),
    .A2(_1588_),
    .ZN(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5578_ (.I(_1618_),
    .Z(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5579_ (.A1(_3303_),
    .A2(_1014_),
    .A3(_1530_),
    .A4(_1589_),
    .ZN(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5580_ (.A1(_3209_),
    .A2(_1118_),
    .ZN(_1621_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5581_ (.A1(_1621_),
    .A2(_1139_),
    .B(_1154_),
    .ZN(_1622_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _5582_ (.A1(_1584_),
    .A2(_1622_),
    .Z(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5583_ (.A1(_1617_),
    .A2(_1619_),
    .B(_1620_),
    .C(_1623_),
    .ZN(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5584_ (.A1(_1614_),
    .A2(_1615_),
    .A3(_1616_),
    .A4(_1624_),
    .ZN(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5585_ (.A1(_1611_),
    .A2(_1625_),
    .ZN(_1626_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5586_ (.A1(_1602_),
    .A2(_1605_),
    .A3(_1626_),
    .ZN(_1627_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5587_ (.A1(_3536_),
    .A2(_0348_),
    .Z(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5588_ (.A1(_3171_),
    .A2(_3173_),
    .A3(_3370_),
    .A4(_3476_),
    .ZN(_1629_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _5589_ (.A1(_3556_),
    .A2(_1628_),
    .A3(_0422_),
    .A4(_1629_),
    .Z(_1630_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _5590_ (.A1(_0480_),
    .A2(_0556_),
    .A3(_0607_),
    .A4(_1630_),
    .ZN(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _5591_ (.A1(_0669_),
    .A2(_1249_),
    .A3(_1436_),
    .A4(_1631_),
    .Z(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5592_ (.A1(_1627_),
    .A2(_1632_),
    .ZN(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5593_ (.I(_1613_),
    .Z(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5594_ (.I(_1563_),
    .Z(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5595_ (.I(_3244_),
    .Z(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5596_ (.I(_1636_),
    .Z(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5597_ (.A1(_1204_),
    .A2(_0657_),
    .ZN(_1638_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5598_ (.I(_1431_),
    .Z(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5599_ (.A1(_1639_),
    .A2(_1156_),
    .B(net49),
    .ZN(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5600_ (.I(_1104_),
    .Z(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5601_ (.A1(net23),
    .A2(_1637_),
    .B1(_1638_),
    .B2(_1640_),
    .C(_1641_),
    .ZN(_1642_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5602_ (.A1(_1121_),
    .A2(_1635_),
    .B(_1642_),
    .ZN(_1643_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5603_ (.A1(_1634_),
    .A2(_1643_),
    .ZN(_1644_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5604_ (.A1(net23),
    .A2(_1633_),
    .ZN(_1645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5605_ (.A1(_1633_),
    .A2(_1644_),
    .B(_1645_),
    .C(_1576_),
    .ZN(_0162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5606_ (.A1(_1317_),
    .A2(_0670_),
    .A3(_1341_),
    .ZN(_1646_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5607_ (.A1(_3149_),
    .A2(_3269_),
    .B(_1421_),
    .ZN(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _5608_ (.A1(_0683_),
    .A2(_0685_),
    .B(_1646_),
    .C(_1647_),
    .ZN(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5609_ (.I(_0682_),
    .Z(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5610_ (.A1(_1146_),
    .A2(_1649_),
    .B(_1609_),
    .ZN(_1650_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5611_ (.I(_1134_),
    .Z(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5612_ (.I(_3207_),
    .Z(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5613_ (.I(_1652_),
    .Z(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5614_ (.A1(_1653_),
    .A2(_1434_),
    .ZN(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5615_ (.A1(_1144_),
    .A2(_1651_),
    .A3(_1525_),
    .A4(_1654_),
    .ZN(_1655_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5616_ (.A1(_1623_),
    .A2(_1648_),
    .A3(_1650_),
    .A4(_1655_),
    .ZN(_1656_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5617_ (.A1(_3316_),
    .A2(_1155_),
    .ZN(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5618_ (.A1(_0863_),
    .A2(_1160_),
    .A3(_1168_),
    .A4(_1657_),
    .ZN(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5619_ (.A1(_1082_),
    .A2(_1321_),
    .A3(_3269_),
    .A4(_0682_),
    .ZN(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5620_ (.A1(_1658_),
    .A2(_1659_),
    .ZN(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5621_ (.A1(_1608_),
    .A2(_1605_),
    .A3(_1656_),
    .A4(_1660_),
    .ZN(_1661_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5622_ (.A1(_1632_),
    .A2(_1661_),
    .ZN(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5623_ (.A1(_1451_),
    .A2(_1517_),
    .ZN(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5624_ (.I(_1489_),
    .Z(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5625_ (.A1(_1555_),
    .A2(_1417_),
    .ZN(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5626_ (.A1(_1417_),
    .A2(_0657_),
    .ZN(_1666_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5627_ (.A1(_1203_),
    .A2(_0674_),
    .ZN(_1667_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5628_ (.A1(_1666_),
    .A2(_1667_),
    .ZN(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5629_ (.A1(_1465_),
    .A2(_1166_),
    .B1(_1665_),
    .B2(_1427_),
    .C(_1668_),
    .ZN(_1669_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5630_ (.A1(_1132_),
    .A2(_1491_),
    .ZN(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5631_ (.A1(net22),
    .A2(_1651_),
    .A3(_1669_),
    .A4(_1670_),
    .ZN(_1671_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5632_ (.A1(_1664_),
    .A2(_1322_),
    .B1(_1345_),
    .B2(_1554_),
    .C(_1671_),
    .ZN(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5633_ (.A1(_1663_),
    .A2(_1672_),
    .ZN(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5634_ (.A1(net22),
    .A2(_1662_),
    .ZN(_1674_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5635_ (.A1(_1662_),
    .A2(_1673_),
    .B(_1674_),
    .C(_1576_),
    .ZN(_0163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5636_ (.I(_1528_),
    .Z(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5637_ (.A1(_3224_),
    .A2(_1495_),
    .A3(_1497_),
    .ZN(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5638_ (.A1(_1675_),
    .A2(_1676_),
    .ZN(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5639_ (.A1(_1618_),
    .A2(_1677_),
    .ZN(_1678_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5640_ (.A1(_1451_),
    .A2(_1317_),
    .ZN(_1679_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5641_ (.A1(_1679_),
    .A2(_1591_),
    .ZN(_1680_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5642_ (.A1(_1523_),
    .A2(_1529_),
    .B(_0862_),
    .ZN(_1681_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5643_ (.A1(_1568_),
    .A2(_1259_),
    .A3(_1680_),
    .A4(_1681_),
    .ZN(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5644_ (.A1(_0862_),
    .A2(_1679_),
    .ZN(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5645_ (.A1(_1420_),
    .A2(_1683_),
    .B(_0919_),
    .ZN(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5646_ (.I(_1519_),
    .Z(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5647_ (.A1(_1685_),
    .A2(_1499_),
    .A3(_1507_),
    .A4(_1599_),
    .ZN(_1686_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _5648_ (.A1(_1678_),
    .A2(_1682_),
    .A3(_1684_),
    .A4(_1686_),
    .ZN(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5649_ (.A1(_3228_),
    .A2(_1634_),
    .B(_1687_),
    .ZN(_1688_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5650_ (.A1(_3186_),
    .A2(_1687_),
    .B(_1688_),
    .C(_1576_),
    .ZN(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5651_ (.I(_1613_),
    .Z(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5652_ (.A1(_3229_),
    .A2(_1689_),
    .B(_1687_),
    .ZN(_1690_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5653_ (.I(_1575_),
    .Z(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5654_ (.A1(_3185_),
    .A2(_1687_),
    .B(_1690_),
    .C(_1691_),
    .ZN(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5655_ (.I(_1266_),
    .Z(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5656_ (.A1(_3311_),
    .A2(_1259_),
    .ZN(_1693_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _5657_ (.A1(_1488_),
    .A2(_1692_),
    .B(_1693_),
    .ZN(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5658_ (.I(_3433_),
    .Z(_1695_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5659_ (.A1(_1695_),
    .A2(_3434_),
    .ZN(_1696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5660_ (.A1(_1153_),
    .A2(_1657_),
    .ZN(_1697_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5661_ (.A1(_0901_),
    .A2(_1138_),
    .ZN(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5662_ (.A1(_1637_),
    .A2(_1698_),
    .B(_1097_),
    .ZN(_1699_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5663_ (.A1(_1696_),
    .A2(_1697_),
    .A3(_1699_),
    .Z(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _5664_ (.I(_1700_),
    .Z(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5665_ (.I0(\as2650.holding_reg[0] ),
    .I1(_1694_),
    .S(_1701_),
    .Z(_1702_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5666_ (.I(_1702_),
    .Z(_0166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5667_ (.I(_1149_),
    .Z(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5668_ (.A1(_1333_),
    .A2(_1703_),
    .ZN(_1704_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5669_ (.I(_1097_),
    .Z(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5670_ (.A1(_3483_),
    .A2(_1705_),
    .ZN(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5671_ (.A1(_1704_),
    .A2(_1706_),
    .ZN(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5672_ (.I0(_3502_),
    .I1(_1707_),
    .S(_1701_),
    .Z(_1708_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5673_ (.I(_1708_),
    .Z(_0167_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5674_ (.A1(_1696_),
    .A2(_1697_),
    .A3(_1699_),
    .ZN(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5675_ (.I(_3528_),
    .Z(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5676_ (.A1(_1241_),
    .A2(_1266_),
    .ZN(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5677_ (.I(_1711_),
    .ZN(_1712_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5678_ (.A1(_1710_),
    .A2(_1641_),
    .B(_1712_),
    .ZN(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5679_ (.A1(_0261_),
    .A2(_1709_),
    .ZN(_1714_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5680_ (.A1(_1709_),
    .A2(_1713_),
    .B(_1714_),
    .ZN(_0168_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5681_ (.I(_1242_),
    .Z(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5682_ (.A1(_1715_),
    .A2(_1105_),
    .ZN(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5683_ (.A1(_0354_),
    .A2(_1705_),
    .ZN(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _5684_ (.A1(_1700_),
    .A2(_1716_),
    .A3(_1717_),
    .Z(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5685_ (.A1(_0281_),
    .A2(_1709_),
    .B(_1718_),
    .ZN(_0169_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5686_ (.I(_1289_),
    .Z(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5687_ (.I(_1719_),
    .Z(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5688_ (.A1(_1720_),
    .A2(_1641_),
    .ZN(_1721_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5689_ (.A1(_0975_),
    .A2(_1705_),
    .ZN(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5690_ (.A1(_1721_),
    .A2(_1722_),
    .ZN(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5691_ (.I0(_0368_),
    .I1(_1723_),
    .S(_1701_),
    .Z(_1724_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5692_ (.I(_1724_),
    .Z(_0170_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5693_ (.A1(_1235_),
    .A2(_1567_),
    .B(_1098_),
    .ZN(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5694_ (.I0(_0458_),
    .I1(_1725_),
    .S(_1701_),
    .Z(_1726_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5695_ (.I(_1726_),
    .Z(_0171_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5696_ (.I(_1700_),
    .Z(_1727_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5697_ (.I(_0547_),
    .Z(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5698_ (.I(_1641_),
    .Z(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5699_ (.A1(_1236_),
    .A2(_1578_),
    .ZN(_1730_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5700_ (.A1(_1728_),
    .A2(_1729_),
    .B(_1730_),
    .ZN(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5701_ (.A1(_0531_),
    .A2(_1727_),
    .ZN(_1732_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5702_ (.A1(_1727_),
    .A2(_1731_),
    .B(_1732_),
    .ZN(_0172_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5703_ (.I(_1259_),
    .Z(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5704_ (.A1(_1554_),
    .A2(_1733_),
    .B(_1267_),
    .ZN(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5705_ (.A1(_1727_),
    .A2(_1734_),
    .ZN(_1735_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5706_ (.A1(_0576_),
    .A2(_1727_),
    .B(_1735_),
    .ZN(_0173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5707_ (.I(_1460_),
    .Z(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5708_ (.A1(_1729_),
    .A2(_1155_),
    .B(_3237_),
    .ZN(_1737_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5709_ (.A1(_1736_),
    .A2(_1737_),
    .Z(_1738_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5710_ (.I(_1738_),
    .Z(_0174_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5711_ (.I(_1568_),
    .Z(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5712_ (.A1(_1739_),
    .A2(_1664_),
    .ZN(_1740_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5713_ (.I(_1204_),
    .Z(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5714_ (.A1(_1439_),
    .A2(_1029_),
    .ZN(_1742_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5715_ (.I(_1742_),
    .Z(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5716_ (.I(_1598_),
    .Z(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5717_ (.I(_1744_),
    .Z(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5718_ (.A1(_1489_),
    .A2(_1426_),
    .ZN(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _5719_ (.A1(_1034_),
    .A2(_1089_),
    .A3(_1066_),
    .A4(_1086_),
    .ZN(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5720_ (.A1(_1745_),
    .A2(_1635_),
    .B1(_1746_),
    .B2(_1747_),
    .ZN(_1748_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5721_ (.I(_1163_),
    .Z(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5722_ (.A1(_1039_),
    .A2(_1749_),
    .A3(_1746_),
    .ZN(_1750_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5723_ (.A1(_1489_),
    .A2(_0685_),
    .B(_1424_),
    .C(_1665_),
    .ZN(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5724_ (.I(_1603_),
    .ZN(_1752_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5725_ (.A1(_1752_),
    .A2(_1631_),
    .ZN(_1753_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5726_ (.A1(_1258_),
    .A2(_1753_),
    .ZN(_1754_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5727_ (.A1(_0662_),
    .A2(_1746_),
    .ZN(_1755_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5728_ (.A1(_1649_),
    .A2(_1754_),
    .A3(_1755_),
    .ZN(_1756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5729_ (.A1(_1751_),
    .A2(_1756_),
    .B(_1427_),
    .ZN(_1757_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5730_ (.A1(_1743_),
    .A2(_1748_),
    .B(_1750_),
    .C(_1757_),
    .ZN(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5731_ (.A1(_1321_),
    .A2(_1345_),
    .B1(_1758_),
    .B2(_1518_),
    .ZN(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5732_ (.A1(_1741_),
    .A2(_1759_),
    .ZN(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5733_ (.A1(_1664_),
    .A2(_3305_),
    .ZN(_1761_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5734_ (.A1(_3184_),
    .A2(_1636_),
    .ZN(_1762_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5735_ (.I(_1500_),
    .Z(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5736_ (.I(_1763_),
    .Z(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5737_ (.A1(_1761_),
    .A2(_1762_),
    .B(_1764_),
    .ZN(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5738_ (.A1(_1527_),
    .A2(_1676_),
    .ZN(_1766_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5739_ (.A1(_1307_),
    .A2(_1636_),
    .B(_1766_),
    .ZN(_1767_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5740_ (.A1(_1555_),
    .A2(_1636_),
    .B(_1763_),
    .ZN(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5741_ (.A1(_1105_),
    .A2(_0687_),
    .A3(_1767_),
    .A4(_1768_),
    .ZN(_1769_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5742_ (.A1(_1578_),
    .A2(_1284_),
    .B1(_1765_),
    .B2(_1769_),
    .C(_1591_),
    .ZN(_1770_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5743_ (.A1(_1586_),
    .A2(_1760_),
    .A3(_1770_),
    .ZN(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5744_ (.I(_1575_),
    .Z(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5745_ (.A1(_1740_),
    .A2(_1771_),
    .B(_1772_),
    .ZN(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5746_ (.I(_1595_),
    .Z(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5747_ (.I(_1577_),
    .Z(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _5748_ (.A1(_0356_),
    .A2(_1752_),
    .A3(_1631_),
    .ZN(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5749_ (.I(_1511_),
    .Z(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5750_ (.A1(_1776_),
    .A2(_1647_),
    .ZN(_1777_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5751_ (.A1(_3149_),
    .A2(_3304_),
    .ZN(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5752_ (.I(_1514_),
    .Z(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5753_ (.I(_1084_),
    .Z(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5754_ (.I(_1780_),
    .Z(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5755_ (.A1(_1781_),
    .A2(_1490_),
    .A3(_1649_),
    .A4(_1778_),
    .ZN(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5756_ (.A1(_1779_),
    .A2(_1782_),
    .ZN(_1783_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5757_ (.A1(_1436_),
    .A2(_1775_),
    .B1(_1777_),
    .B2(_1778_),
    .C(_1783_),
    .ZN(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5758_ (.I(_1695_),
    .Z(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5759_ (.I(_1530_),
    .Z(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5760_ (.I(_1786_),
    .Z(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5761_ (.A1(_1778_),
    .A2(_1762_),
    .A3(_1768_),
    .ZN(_1788_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5762_ (.A1(_1149_),
    .A2(_1490_),
    .A3(_1767_),
    .ZN(_1789_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5763_ (.A1(_1787_),
    .A2(_1788_),
    .B(_1789_),
    .ZN(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5764_ (.A1(_1096_),
    .A2(_1747_),
    .ZN(_1791_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5765_ (.A1(_1030_),
    .A2(_1039_),
    .B1(_1778_),
    .B2(_1781_),
    .C(_1078_),
    .ZN(_1792_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5766_ (.A1(_1791_),
    .A2(_1792_),
    .ZN(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5767_ (.A1(_1785_),
    .A2(_1441_),
    .A3(_1790_),
    .B(_1793_),
    .ZN(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5768_ (.A1(_1774_),
    .A2(_1784_),
    .A3(_1794_),
    .ZN(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5769_ (.A1(_1739_),
    .A2(_1082_),
    .B(_1795_),
    .ZN(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5770_ (.A1(_1773_),
    .A2(_1796_),
    .ZN(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5771_ (.I(_1774_),
    .Z(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5772_ (.I(_1575_),
    .Z(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5773_ (.A1(_1143_),
    .A2(_1589_),
    .ZN(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5774_ (.I(_1799_),
    .Z(_1800_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5775_ (.I(_1800_),
    .Z(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5776_ (.I(_1423_),
    .Z(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5777_ (.A1(_0655_),
    .A2(_3219_),
    .Z(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5778_ (.A1(_1664_),
    .A2(_3269_),
    .B(_1803_),
    .ZN(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5779_ (.A1(_1802_),
    .A2(_1665_),
    .A3(_1804_),
    .ZN(_1805_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5780_ (.I(_0663_),
    .Z(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5781_ (.I(_1806_),
    .Z(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5782_ (.A1(_1807_),
    .A2(_1803_),
    .ZN(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5783_ (.A1(_1639_),
    .A2(_1808_),
    .B(_1327_),
    .C(_0654_),
    .ZN(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5784_ (.A1(_1153_),
    .A2(_1803_),
    .Z(_1810_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5785_ (.I(_1325_),
    .Z(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5786_ (.I(_1811_),
    .Z(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5787_ (.A1(_1805_),
    .A2(_1809_),
    .B1(_1810_),
    .B2(_1812_),
    .ZN(_1813_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5788_ (.A1(_1651_),
    .A2(_1090_),
    .B(_1803_),
    .ZN(_1814_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5789_ (.I(_1494_),
    .Z(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5790_ (.A1(_1815_),
    .A2(_1635_),
    .ZN(_1816_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5791_ (.A1(_1814_),
    .A2(_1816_),
    .Z(_1817_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5792_ (.I(_1029_),
    .Z(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5793_ (.A1(_3220_),
    .A2(_1818_),
    .B(_1463_),
    .ZN(_1819_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5794_ (.A1(_1466_),
    .A2(_1813_),
    .B1(_1817_),
    .B2(_1819_),
    .ZN(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5795_ (.A1(_3251_),
    .A2(_1657_),
    .A3(_1698_),
    .B(_1808_),
    .ZN(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5796_ (.A1(_1801_),
    .A2(_1820_),
    .B1(_1821_),
    .B2(_1619_),
    .C(_1774_),
    .ZN(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5797_ (.A1(_1797_),
    .A2(_0655_),
    .B(_1798_),
    .C(_1822_),
    .ZN(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5798_ (.A1(_3215_),
    .A2(_3217_),
    .A3(_3360_),
    .ZN(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5799_ (.A1(_0655_),
    .A2(_3219_),
    .B(_3268_),
    .ZN(_1824_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5800_ (.A1(_1823_),
    .A2(_1824_),
    .ZN(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5801_ (.A1(_1572_),
    .A2(_1825_),
    .ZN(_1826_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5802_ (.A1(_0674_),
    .A2(_1666_),
    .B(_1826_),
    .ZN(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5803_ (.I(_1766_),
    .Z(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5804_ (.A1(_3314_),
    .A2(_1828_),
    .B(_1637_),
    .ZN(_1829_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5805_ (.A1(_1762_),
    .A2(_1825_),
    .A3(_1829_),
    .ZN(_1830_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5806_ (.I(_1766_),
    .Z(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5807_ (.I(_1831_),
    .Z(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5808_ (.A1(_1553_),
    .A2(_1637_),
    .ZN(_1833_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5809_ (.I(_1695_),
    .Z(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5810_ (.A1(_1832_),
    .A2(_1833_),
    .B(_1834_),
    .C(_0657_),
    .ZN(_1835_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5811_ (.A1(_1554_),
    .A2(_1153_),
    .A3(_1776_),
    .B(_1454_),
    .ZN(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5812_ (.I(_1779_),
    .Z(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5813_ (.A1(_1830_),
    .A2(_1835_),
    .B1(_1836_),
    .B2(_1837_),
    .C(_1577_),
    .ZN(_1838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5814_ (.A1(_1797_),
    .A2(_3268_),
    .B1(_1827_),
    .B2(_1838_),
    .C(_1798_),
    .ZN(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5815_ (.I(\as2650.cycle[4] ),
    .Z(_1839_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5816_ (.A1(_1568_),
    .A2(_1823_),
    .ZN(_1840_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5817_ (.A1(_1839_),
    .A2(_1840_),
    .B(_1470_),
    .ZN(_1841_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5818_ (.A1(_1839_),
    .A2(_1840_),
    .B(_1841_),
    .ZN(_0179_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5819_ (.A1(_1839_),
    .A2(_1840_),
    .ZN(_1842_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5820_ (.A1(\as2650.cycle[5] ),
    .A2(_1842_),
    .Z(_1843_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5821_ (.A1(_1773_),
    .A2(_1843_),
    .ZN(_0180_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5822_ (.A1(\as2650.cycle[5] ),
    .A2(_1839_),
    .ZN(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5823_ (.A1(_1675_),
    .A2(_1823_),
    .A3(_1844_),
    .Z(_1845_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5824_ (.A1(_1823_),
    .A2(_1844_),
    .B(_1675_),
    .ZN(_1846_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5825_ (.I(_1831_),
    .Z(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5826_ (.A1(_3184_),
    .A2(_3314_),
    .A3(_1847_),
    .B(_1619_),
    .ZN(_1848_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5827_ (.A1(_1845_),
    .A2(_1846_),
    .A3(_1848_),
    .ZN(_1849_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5828_ (.I(_1250_),
    .Z(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5829_ (.A1(_1654_),
    .A2(_1850_),
    .ZN(_1851_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5830_ (.A1(_1739_),
    .A2(_1620_),
    .A3(_1851_),
    .ZN(_1852_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5831_ (.I(_1115_),
    .Z(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5832_ (.A1(_1739_),
    .A2(_1675_),
    .B1(_1849_),
    .B2(_1852_),
    .C(_1853_),
    .ZN(_0181_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5833_ (.I(_1162_),
    .Z(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5834_ (.I(_1854_),
    .Z(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _5835_ (.A1(_1733_),
    .A2(_1764_),
    .A3(_1847_),
    .B(_1619_),
    .ZN(_1856_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5836_ (.A1(_3141_),
    .A2(_1845_),
    .Z(_1857_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5837_ (.A1(_1855_),
    .A2(_1590_),
    .B1(_1856_),
    .B2(_1857_),
    .C(_1774_),
    .ZN(_1858_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5838_ (.A1(_1797_),
    .A2(_3141_),
    .B(_1798_),
    .C(_1858_),
    .ZN(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5839_ (.A1(_1578_),
    .A2(_1071_),
    .B1(_1178_),
    .B2(_1061_),
    .C(net9),
    .ZN(_1859_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5840_ (.A1(_1130_),
    .A2(_1351_),
    .ZN(_1860_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5841_ (.A1(_1295_),
    .A2(_1351_),
    .B(_1860_),
    .ZN(_1861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5842_ (.A1(_1071_),
    .A2(_1267_),
    .B(_3237_),
    .ZN(_1862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5843_ (.A1(_1179_),
    .A2(_1861_),
    .B(_1862_),
    .ZN(_1863_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5844_ (.A1(_1295_),
    .A2(_1797_),
    .B1(_1859_),
    .B2(_1863_),
    .C(_1853_),
    .ZN(_0183_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5845_ (.A1(_1609_),
    .A2(_1610_),
    .ZN(_1864_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5846_ (.A1(_1621_),
    .A2(_1139_),
    .ZN(_1865_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5847_ (.A1(_1059_),
    .A2(_1064_),
    .B(_1865_),
    .ZN(_1866_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _5848_ (.A1(_1517_),
    .A2(_1579_),
    .B1(_1866_),
    .B2(_1032_),
    .C(_1663_),
    .ZN(_1867_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5849_ (.A1(_1607_),
    .A2(_1864_),
    .A3(_1867_),
    .ZN(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5850_ (.A1(_1517_),
    .A2(_1163_),
    .ZN(_1869_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5851_ (.A1(_1442_),
    .A2(_1600_),
    .ZN(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5852_ (.A1(_0357_),
    .A2(_1869_),
    .B(_1870_),
    .ZN(_1871_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5853_ (.A1(_1014_),
    .A2(_1523_),
    .A3(_1341_),
    .ZN(_1872_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5854_ (.A1(_0868_),
    .A2(_1064_),
    .ZN(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5855_ (.A1(_1174_),
    .A2(_1873_),
    .B(_1032_),
    .ZN(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5856_ (.A1(_1681_),
    .A2(_1872_),
    .A3(_1874_),
    .ZN(_1875_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5857_ (.A1(_0659_),
    .A2(_1416_),
    .A3(_1422_),
    .ZN(_1876_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _5858_ (.A1(_3271_),
    .A2(_1420_),
    .A3(_1422_),
    .A4(_1646_),
    .ZN(_1877_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5859_ (.A1(_1648_),
    .A2(_1877_),
    .ZN(_1878_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5860_ (.A1(_1684_),
    .A2(_1875_),
    .A3(_1876_),
    .A4(_1878_),
    .ZN(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5861_ (.A1(_3433_),
    .A2(_1456_),
    .B(_1879_),
    .ZN(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5862_ (.A1(_1660_),
    .A2(_1868_),
    .A3(_1871_),
    .A4(_1880_),
    .ZN(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5863_ (.I(_1881_),
    .Z(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5864_ (.I(_1882_),
    .Z(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5865_ (.A1(_0864_),
    .A2(_1613_),
    .ZN(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5866_ (.I(_1884_),
    .Z(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5867_ (.I(_1881_),
    .Z(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5868_ (.A1(_0646_),
    .A2(_1885_),
    .B(_1886_),
    .ZN(_1887_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5869_ (.A1(_1426_),
    .A2(_1423_),
    .B(_1775_),
    .ZN(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5870_ (.I(_1888_),
    .Z(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5871_ (.I(_1055_),
    .Z(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5872_ (.I(\as2650.addr_buff[0] ),
    .Z(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5873_ (.A1(_1891_),
    .A2(_1562_),
    .ZN(_1892_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5874_ (.I(_0664_),
    .Z(_1893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5875_ (.A1(_3374_),
    .A2(_1893_),
    .ZN(_1894_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _5876_ (.A1(_1890_),
    .A2(_1892_),
    .A3(_1894_),
    .ZN(_1895_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5877_ (.A1(_0643_),
    .A2(_3373_),
    .Z(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5878_ (.I(_0643_),
    .Z(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5879_ (.I(_1324_),
    .Z(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5880_ (.A1(_1897_),
    .A2(_1898_),
    .ZN(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5881_ (.A1(_1433_),
    .A2(_1896_),
    .B(_1899_),
    .C(_1435_),
    .ZN(_1900_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5882_ (.A1(_1431_),
    .A2(_1900_),
    .ZN(_1901_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5883_ (.A1(_1488_),
    .A2(_3293_),
    .Z(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5884_ (.A1(_3374_),
    .A2(_0664_),
    .ZN(_1903_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5885_ (.A1(_1893_),
    .A2(_1902_),
    .B(_1903_),
    .C(_1509_),
    .ZN(_1904_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5886_ (.A1(_1895_),
    .A2(_1901_),
    .B(_1904_),
    .ZN(_1905_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5887_ (.A1(_1149_),
    .A2(_1905_),
    .ZN(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5888_ (.A1(_0645_),
    .A2(_1338_),
    .ZN(_1907_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5889_ (.A1(_1154_),
    .A2(_1753_),
    .ZN(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5890_ (.I(_1908_),
    .Z(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _5891_ (.A1(_1639_),
    .A2(_1899_),
    .A3(_1907_),
    .A4(_1909_),
    .ZN(_1910_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5892_ (.A1(_0645_),
    .A2(_1889_),
    .B(_1906_),
    .C(_1910_),
    .ZN(_1911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5893_ (.A1(_1034_),
    .A2(_1511_),
    .ZN(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5894_ (.A1(_1033_),
    .A2(_1325_),
    .ZN(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5895_ (.I(_1913_),
    .Z(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5896_ (.I(_1914_),
    .Z(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5897_ (.A1(_1896_),
    .A2(_1915_),
    .B(_1463_),
    .ZN(_1916_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5898_ (.A1(_1345_),
    .A2(_1911_),
    .B1(_1912_),
    .B2(_1897_),
    .C(_1916_),
    .ZN(_1917_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5899_ (.I(_1151_),
    .Z(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5900_ (.A1(_1142_),
    .A2(_1096_),
    .ZN(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5901_ (.A1(\as2650.stack_ptr[2] ),
    .A2(_0648_),
    .ZN(_1920_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5902_ (.I(_1920_),
    .Z(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5903_ (.I(_1921_),
    .Z(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5904_ (.A1(\as2650.stack[1][0] ),
    .A2(_0782_),
    .B1(_0806_),
    .B2(\as2650.stack[0][0] ),
    .ZN(_1923_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5905_ (.I(_0752_),
    .Z(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5906_ (.I(_1924_),
    .Z(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5907_ (.A1(_0652_),
    .A2(\as2650.stack[3][0] ),
    .B1(\as2650.stack[2][0] ),
    .B2(_1925_),
    .ZN(_1926_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5908_ (.A1(_1922_),
    .A2(_1923_),
    .A3(_1926_),
    .ZN(_1927_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5909_ (.A1(\as2650.stack[5][0] ),
    .A2(_0782_),
    .B1(_0806_),
    .B2(\as2650.stack[4][0] ),
    .ZN(_1928_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5910_ (.I(_0649_),
    .Z(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5911_ (.A1(\as2650.stack[7][0] ),
    .A2(_1929_),
    .B1(_1925_),
    .B2(\as2650.stack[6][0] ),
    .ZN(_1930_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5912_ (.A1(_1473_),
    .A2(_1928_),
    .A3(_1930_),
    .ZN(_1931_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _5913_ (.A1(_1919_),
    .A2(_1927_),
    .A3(_1931_),
    .ZN(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5914_ (.A1(_1897_),
    .A2(_1918_),
    .B(_1932_),
    .ZN(_1933_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5915_ (.A1(_1917_),
    .A2(_1933_),
    .B(_1801_),
    .ZN(_1934_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5916_ (.A1(_0646_),
    .A2(_1883_),
    .B1(_1887_),
    .B2(_1934_),
    .C(_1853_),
    .ZN(_0184_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5917_ (.I(_1882_),
    .Z(_1935_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5918_ (.I(_1935_),
    .Z(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5919_ (.I(\as2650.pc[1] ),
    .Z(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5920_ (.A1(_1937_),
    .A2(_0643_),
    .Z(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5921_ (.I(_1884_),
    .Z(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5922_ (.A1(_1067_),
    .A2(_1326_),
    .ZN(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5923_ (.A1(_0695_),
    .A2(_0642_),
    .Z(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5924_ (.A1(_0642_),
    .A2(_3155_),
    .ZN(_1942_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5925_ (.A1(_0695_),
    .A2(_1942_),
    .Z(_1943_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5926_ (.A1(_3466_),
    .A2(_1512_),
    .ZN(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5927_ (.A1(\as2650.addr_buff[1] ),
    .A2(_1127_),
    .B(_1422_),
    .C(_1054_),
    .ZN(_1945_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5928_ (.A1(\as2650.pc[0] ),
    .A2(net1),
    .ZN(_1946_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5929_ (.A1(\as2650.pc[1] ),
    .A2(net2),
    .ZN(_1947_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5930_ (.A1(_1946_),
    .A2(_1947_),
    .Z(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5931_ (.A1(_1336_),
    .A2(_1948_),
    .ZN(_1949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5932_ (.A1(_1337_),
    .A2(_1941_),
    .B(_1949_),
    .ZN(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5933_ (.A1(_1133_),
    .A2(_1950_),
    .B(_1124_),
    .ZN(_1951_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5934_ (.A1(_1944_),
    .A2(_1945_),
    .B1(_1951_),
    .B2(_1430_),
    .ZN(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5935_ (.A1(_1775_),
    .A2(_1938_),
    .B1(_1943_),
    .B2(_1908_),
    .C(_1952_),
    .ZN(_1953_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5936_ (.A1(_1157_),
    .A2(_1941_),
    .ZN(_1954_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5937_ (.A1(net1),
    .A2(_3293_),
    .Z(_1955_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5938_ (.I0(\as2650.r123[2][1] ),
    .I1(\as2650.r123_2[2][1] ),
    .S(_3324_),
    .Z(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5939_ (.A1(net2),
    .A2(_1956_),
    .Z(_1957_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _5940_ (.A1(_1955_),
    .A2(_1957_),
    .ZN(_1958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5941_ (.A1(_3465_),
    .A2(_1127_),
    .ZN(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5942_ (.A1(_1598_),
    .A2(_1958_),
    .B(_1959_),
    .C(_1145_),
    .ZN(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5943_ (.A1(_1249_),
    .A2(_1938_),
    .B1(_1954_),
    .B2(_1960_),
    .C(_0682_),
    .ZN(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _5944_ (.A1(_1326_),
    .A2(_1953_),
    .A3(_1961_),
    .Z(_1962_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _5945_ (.A1(_1067_),
    .A2(_1343_),
    .ZN(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5946_ (.A1(_1963_),
    .A2(_1948_),
    .ZN(_1964_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _5947_ (.A1(_1940_),
    .A2(_1941_),
    .B(_1962_),
    .C(_1964_),
    .ZN(_1965_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5948_ (.I(_1142_),
    .Z(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5949_ (.I(_0648_),
    .Z(_1967_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5950_ (.I(_1967_),
    .Z(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5951_ (.I(_0753_),
    .Z(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5952_ (.I(_0780_),
    .Z(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5953_ (.I(_0804_),
    .Z(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5954_ (.A1(\as2650.stack[1][1] ),
    .A2(_1970_),
    .B1(_1971_),
    .B2(\as2650.stack[0][1] ),
    .ZN(_1972_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5955_ (.I(_1972_),
    .ZN(_1973_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5956_ (.A1(\as2650.stack[3][1] ),
    .A2(_1968_),
    .B1(_1969_),
    .B2(\as2650.stack[2][1] ),
    .C(_1973_),
    .ZN(_1974_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5957_ (.I(_1970_),
    .Z(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5958_ (.I(_1971_),
    .Z(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5959_ (.I(_0753_),
    .Z(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _5960_ (.A1(\as2650.stack[5][1] ),
    .A2(_1975_),
    .B1(_1976_),
    .B2(\as2650.stack[4][1] ),
    .C1(\as2650.stack[6][1] ),
    .C2(_1977_),
    .ZN(_1978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5961_ (.A1(\as2650.stack[7][1] ),
    .A2(_0650_),
    .B(_1921_),
    .ZN(_1979_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5962_ (.A1(_1922_),
    .A2(_1974_),
    .B1(_1978_),
    .B2(_1979_),
    .C(_1749_),
    .ZN(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _5963_ (.A1(_1743_),
    .A2(_1938_),
    .B1(_1965_),
    .B2(_1966_),
    .C(_1980_),
    .ZN(_1981_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5964_ (.A1(_1939_),
    .A2(_1981_),
    .ZN(_1982_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5965_ (.A1(_1885_),
    .A2(_1938_),
    .B(_1982_),
    .C(_1886_),
    .ZN(_1983_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _5966_ (.A1(_0696_),
    .A2(_1936_),
    .B(_1983_),
    .C(_1691_),
    .ZN(_0185_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5967_ (.I(_1935_),
    .Z(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5968_ (.I(_1882_),
    .Z(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _5969_ (.A1(\as2650.pc[2] ),
    .A2(_1937_),
    .A3(\as2650.pc[0] ),
    .ZN(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5970_ (.A1(_0696_),
    .A2(_0644_),
    .B(_0699_),
    .ZN(_1987_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _5971_ (.A1(_1986_),
    .A2(_1987_),
    .ZN(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5972_ (.I(_1889_),
    .Z(_1989_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5973_ (.I(_1940_),
    .Z(_1990_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5974_ (.A1(_0699_),
    .A2(_1239_),
    .Z(_1991_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5975_ (.A1(\as2650.pc[1] ),
    .A2(_3462_),
    .ZN(_1992_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5976_ (.A1(_1946_),
    .A2(_1947_),
    .B(_1992_),
    .ZN(_1993_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5977_ (.A1(_1991_),
    .A2(_1993_),
    .Z(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _5978_ (.I(_1439_),
    .Z(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _5979_ (.A1(_1990_),
    .A2(_1988_),
    .B1(_1994_),
    .B2(_1915_),
    .C(_1995_),
    .ZN(_1996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5980_ (.I(_1799_),
    .Z(_1997_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5981_ (.A1(_1989_),
    .A2(_1996_),
    .B(_1997_),
    .ZN(_1998_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5982_ (.I(_1327_),
    .Z(_1999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5983_ (.I(_1525_),
    .Z(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5984_ (.A1(_0695_),
    .A2(_1942_),
    .ZN(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _5985_ (.A1(_0700_),
    .A2(_2001_),
    .Z(_2002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _5986_ (.I(\as2650.addr_buff[2] ),
    .ZN(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5987_ (.I(_1452_),
    .Z(_2004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _5988_ (.A1(_1240_),
    .A2(_2004_),
    .ZN(_2005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5989_ (.A1(_2003_),
    .A2(_2004_),
    .B(_2005_),
    .ZN(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5990_ (.I(_1337_),
    .Z(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _5991_ (.A1(_2007_),
    .A2(_1988_),
    .B(_1055_),
    .ZN(_2008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _5992_ (.I(_1324_),
    .Z(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _5993_ (.A1(_2009_),
    .A2(_1994_),
    .ZN(_2010_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _5994_ (.A1(_1890_),
    .A2(_2006_),
    .B1(_2008_),
    .B2(_2010_),
    .ZN(_2011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _5995_ (.A1(_1909_),
    .A2(_2002_),
    .B1(_2011_),
    .B2(_1104_),
    .ZN(_2012_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _5996_ (.I(_1893_),
    .Z(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _5997_ (.I0(\as2650.r123[2][2] ),
    .I1(\as2650.r123_2[2][2] ),
    .S(_3194_),
    .Z(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _5998_ (.A1(_3462_),
    .A2(_1956_),
    .Z(_2015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _5999_ (.A1(_1955_),
    .A2(_1957_),
    .B(_2015_),
    .ZN(_2016_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6000_ (.A1(_1239_),
    .A2(_2014_),
    .A3(_2016_),
    .Z(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6001_ (.A1(_1240_),
    .A2(_0664_),
    .ZN(_2018_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6002_ (.A1(_1157_),
    .A2(_1430_),
    .ZN(_2019_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6003_ (.I(_2019_),
    .Z(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6004_ (.A1(_2013_),
    .A2(_2017_),
    .B(_2018_),
    .C(_2020_),
    .ZN(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6005_ (.A1(_2000_),
    .A2(_2012_),
    .B(_2021_),
    .ZN(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6006_ (.A1(_1999_),
    .A2(_2022_),
    .ZN(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6007_ (.I(_1472_),
    .Z(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6008_ (.I(_1970_),
    .Z(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6009_ (.A1(\as2650.stack[6][2] ),
    .A2(_1969_),
    .B1(_2025_),
    .B2(\as2650.stack[5][2] ),
    .ZN(_2026_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6010_ (.I(_1971_),
    .Z(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6011_ (.A1(\as2650.stack[7][2] ),
    .A2(_1968_),
    .B1(_2027_),
    .B2(\as2650.stack[4][2] ),
    .ZN(_2028_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6012_ (.A1(_2024_),
    .A2(_2026_),
    .A3(_2028_),
    .ZN(_2029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6013_ (.I(_1920_),
    .Z(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6014_ (.A1(\as2650.stack[3][2] ),
    .A2(_1968_),
    .B1(_1977_),
    .B2(\as2650.stack[2][2] ),
    .ZN(_2031_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6015_ (.A1(\as2650.stack[1][2] ),
    .A2(_2025_),
    .B1(_1976_),
    .B2(\as2650.stack[0][2] ),
    .ZN(_2032_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6016_ (.A1(_2030_),
    .A2(_2031_),
    .A3(_2032_),
    .ZN(_2033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6017_ (.A1(_2029_),
    .A2(_2033_),
    .ZN(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6018_ (.A1(_1743_),
    .A2(_1988_),
    .B1(_2034_),
    .B2(_1919_),
    .ZN(_2035_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6019_ (.A1(_1996_),
    .A2(_2023_),
    .B(_2035_),
    .ZN(_2036_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6020_ (.I(_1800_),
    .Z(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6021_ (.A1(_1988_),
    .A2(_1998_),
    .B1(_2036_),
    .B2(_2037_),
    .ZN(_2038_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6022_ (.I(_1469_),
    .Z(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6023_ (.A1(_1985_),
    .A2(_2038_),
    .B(_2039_),
    .ZN(_2040_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6024_ (.A1(_0702_),
    .A2(_1984_),
    .B(_2040_),
    .ZN(_0186_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6025_ (.I(\as2650.pc[3] ),
    .Z(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6026_ (.A1(_2041_),
    .A2(_1986_),
    .Z(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6027_ (.A1(\as2650.pc[3] ),
    .A2(net4),
    .ZN(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6028_ (.A1(_0704_),
    .A2(_1297_),
    .ZN(_2044_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6029_ (.A1(_2043_),
    .A2(_2044_),
    .ZN(_2045_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6030_ (.A1(\as2650.pc[2] ),
    .A2(net3),
    .Z(_2046_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6031_ (.A1(_0699_),
    .A2(_3539_),
    .ZN(_2047_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6032_ (.A1(_2046_),
    .A2(_1993_),
    .B(_2047_),
    .ZN(_2048_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6033_ (.A1(_2045_),
    .A2(_2048_),
    .ZN(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6034_ (.A1(_1963_),
    .A2(_2049_),
    .ZN(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6035_ (.A1(_1990_),
    .A2(_2042_),
    .B(_2050_),
    .C(_1966_),
    .ZN(_2051_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6036_ (.A1(_1989_),
    .A2(_2051_),
    .B(_1997_),
    .ZN(_2052_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6037_ (.A1(_1084_),
    .A2(_1423_),
    .ZN(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6038_ (.I(_2053_),
    .Z(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6039_ (.A1(_1715_),
    .A2(_1745_),
    .B(_2054_),
    .ZN(_2055_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6040_ (.I(_1453_),
    .Z(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6041_ (.A1(_3538_),
    .A2(_2014_),
    .ZN(_2057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6042_ (.A1(_3538_),
    .A2(_2014_),
    .ZN(_2058_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6043_ (.A1(_2016_),
    .A2(_2057_),
    .B(_2058_),
    .ZN(_2059_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6044_ (.I0(\as2650.r123[2][3] ),
    .I1(\as2650.r123_2[2][3] ),
    .S(_3325_),
    .Z(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6045_ (.A1(_0343_),
    .A2(_2060_),
    .Z(_2061_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6046_ (.A1(_2059_),
    .A2(_2061_),
    .Z(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6047_ (.A1(_2056_),
    .A2(_2062_),
    .ZN(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6048_ (.I(_1811_),
    .Z(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6049_ (.I(_1525_),
    .Z(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6050_ (.I(_1908_),
    .Z(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6051_ (.A1(\as2650.pc[2] ),
    .A2(_2001_),
    .ZN(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6052_ (.A1(_2041_),
    .A2(_2067_),
    .Z(_2068_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6053_ (.A1(_2009_),
    .A2(_2042_),
    .ZN(_2069_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6054_ (.A1(_1653_),
    .A2(_2049_),
    .B(_2069_),
    .C(_1435_),
    .ZN(_2070_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6055_ (.A1(_1242_),
    .A2(_1513_),
    .B1(_1815_),
    .B2(\as2650.addr_buff[3] ),
    .C(_1210_),
    .ZN(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6056_ (.A1(_2066_),
    .A2(_2068_),
    .B1(_2070_),
    .B2(_2071_),
    .ZN(_2072_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6057_ (.A1(_2065_),
    .A2(_2072_),
    .ZN(_2073_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6058_ (.A1(_2055_),
    .A2(_2063_),
    .B(_2064_),
    .C(_2073_),
    .ZN(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6059_ (.I(_1967_),
    .Z(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6060_ (.I(_0780_),
    .Z(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6061_ (.A1(\as2650.stack[7][3] ),
    .A2(_2075_),
    .B1(_2076_),
    .B2(\as2650.stack[5][3] ),
    .ZN(_2077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6062_ (.I(_0753_),
    .Z(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6063_ (.I(_0804_),
    .Z(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6064_ (.A1(\as2650.stack[6][3] ),
    .A2(_2078_),
    .B1(_2079_),
    .B2(\as2650.stack[4][3] ),
    .ZN(_2080_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6065_ (.A1(_2024_),
    .A2(_2077_),
    .A3(_2080_),
    .ZN(_2081_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6066_ (.I(_0780_),
    .Z(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6067_ (.A1(\as2650.stack[3][3] ),
    .A2(_2075_),
    .B1(_2082_),
    .B2(\as2650.stack[1][3] ),
    .ZN(_2083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6068_ (.I(_0804_),
    .Z(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6069_ (.A1(\as2650.stack[2][3] ),
    .A2(_2078_),
    .B1(_2084_),
    .B2(\as2650.stack[0][3] ),
    .ZN(_2085_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6070_ (.A1(_2030_),
    .A2(_2083_),
    .A3(_2085_),
    .ZN(_2086_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6071_ (.A1(_1030_),
    .A2(_2081_),
    .A3(_2086_),
    .ZN(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6072_ (.I(_1455_),
    .Z(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6073_ (.A1(_1818_),
    .A2(_2042_),
    .B(_2087_),
    .C(_2088_),
    .ZN(_2089_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6074_ (.A1(_2051_),
    .A2(_2074_),
    .B(_2089_),
    .ZN(_2090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6075_ (.A1(_2042_),
    .A2(_2052_),
    .B1(_2090_),
    .B2(_2037_),
    .ZN(_2091_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6076_ (.A1(_1985_),
    .A2(_2091_),
    .B(_2039_),
    .ZN(_2092_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6077_ (.A1(_0706_),
    .A2(_1984_),
    .B(_2092_),
    .ZN(_0187_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6078_ (.A1(_0705_),
    .A2(_1986_),
    .ZN(_2093_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6079_ (.A1(_0709_),
    .A2(_2093_),
    .Z(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6080_ (.I(_1940_),
    .Z(_2095_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6081_ (.A1(_0708_),
    .A2(net5),
    .Z(_2096_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6082_ (.I(_2096_),
    .ZN(_2097_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6083_ (.A1(_2046_),
    .A2(_1993_),
    .B(_2044_),
    .C(_2047_),
    .ZN(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6084_ (.A1(_2043_),
    .A2(_2098_),
    .Z(_2099_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6085_ (.A1(_2097_),
    .A2(_2099_),
    .Z(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _6086_ (.I(_1914_),
    .Z(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6087_ (.A1(_2095_),
    .A2(_2094_),
    .B1(_2100_),
    .B2(_2101_),
    .C(_1995_),
    .ZN(_2102_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6088_ (.A1(_1989_),
    .A2(_2102_),
    .B(_1997_),
    .ZN(_2103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6089_ (.A1(_0704_),
    .A2(_2067_),
    .ZN(_2104_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6090_ (.A1(_0709_),
    .A2(_2104_),
    .Z(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6091_ (.A1(_1337_),
    .A2(_2094_),
    .Z(_2106_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6092_ (.A1(_1898_),
    .A2(_2100_),
    .B(_2106_),
    .C(_3222_),
    .ZN(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6093_ (.A1(_1719_),
    .A2(_1893_),
    .B1(_1128_),
    .B2(\as2650.addr_buff[4] ),
    .C(_2107_),
    .ZN(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6094_ (.A1(_1909_),
    .A2(_2105_),
    .B1(_2108_),
    .B2(_1104_),
    .ZN(_2109_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6095_ (.I0(\as2650.r123[2][4] ),
    .I1(\as2650.r123_2[2][4] ),
    .S(_3194_),
    .Z(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6096_ (.A1(_0343_),
    .A2(_2060_),
    .Z(_2111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6097_ (.A1(_2059_),
    .A2(_2061_),
    .B(_2111_),
    .ZN(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6098_ (.A1(_1289_),
    .A2(_2110_),
    .A3(_2112_),
    .Z(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6099_ (.A1(_1289_),
    .A2(_1806_),
    .ZN(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6100_ (.A1(_2013_),
    .A2(_2113_),
    .B(_2114_),
    .C(_2020_),
    .ZN(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6101_ (.A1(_2000_),
    .A2(_2109_),
    .B(_2115_),
    .ZN(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6102_ (.A1(_1999_),
    .A2(_2116_),
    .ZN(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6103_ (.A1(\as2650.stack[7][4] ),
    .A2(_2075_),
    .B1(_2076_),
    .B2(\as2650.stack[5][4] ),
    .ZN(_2118_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6104_ (.A1(\as2650.stack[6][4] ),
    .A2(_2078_),
    .B1(_2079_),
    .B2(\as2650.stack[4][4] ),
    .ZN(_2119_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6105_ (.A1(_2024_),
    .A2(_2118_),
    .A3(_2119_),
    .ZN(_2120_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6106_ (.A1(\as2650.stack[3][4] ),
    .A2(_2075_),
    .B1(_2082_),
    .B2(\as2650.stack[1][4] ),
    .ZN(_2121_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6107_ (.I(_0752_),
    .Z(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6108_ (.A1(\as2650.stack[2][4] ),
    .A2(_2122_),
    .B1(_2084_),
    .B2(\as2650.stack[0][4] ),
    .ZN(_2123_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6109_ (.A1(_1921_),
    .A2(_2121_),
    .A3(_2123_),
    .ZN(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6110_ (.A1(_1030_),
    .A2(_2120_),
    .A3(_2124_),
    .ZN(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6111_ (.A1(_1818_),
    .A2(_2094_),
    .B(_2125_),
    .C(_2088_),
    .ZN(_2126_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6112_ (.A1(_2102_),
    .A2(_2117_),
    .B(_2126_),
    .ZN(_2127_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6113_ (.A1(_2094_),
    .A2(_2103_),
    .B1(_2127_),
    .B2(_2037_),
    .ZN(_2128_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6114_ (.A1(_1985_),
    .A2(_2128_),
    .B(_2039_),
    .ZN(_2129_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6115_ (.A1(_0711_),
    .A2(_1984_),
    .B(_2129_),
    .ZN(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6116_ (.I(_1882_),
    .Z(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6117_ (.A1(_0709_),
    .A2(_0704_),
    .A3(_1986_),
    .ZN(_2131_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6118_ (.A1(_0716_),
    .A2(_2131_),
    .Z(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6119_ (.A1(\as2650.pc[5] ),
    .A2(net6),
    .ZN(_2133_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6120_ (.I(_2133_),
    .ZN(_2134_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6121_ (.I(\as2650.pc[4] ),
    .Z(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6122_ (.A1(_2096_),
    .A2(_2099_),
    .ZN(_2136_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6123_ (.A1(_2135_),
    .A2(_1270_),
    .B(_2136_),
    .ZN(_2137_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6124_ (.A1(_2134_),
    .A2(_2137_),
    .Z(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6125_ (.A1(_2095_),
    .A2(_2132_),
    .B1(_2138_),
    .B2(_2101_),
    .C(_1995_),
    .ZN(_2139_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6126_ (.A1(_1989_),
    .A2(_2139_),
    .B(_1997_),
    .ZN(_2140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6127_ (.I(_0715_),
    .Z(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6128_ (.A1(_2141_),
    .A2(\as2650.pc[4] ),
    .A3(_2104_),
    .ZN(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6129_ (.A1(_2135_),
    .A2(_2104_),
    .ZN(_2143_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6130_ (.A1(_0717_),
    .A2(_2143_),
    .ZN(_2144_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6131_ (.A1(_2142_),
    .A2(_2144_),
    .ZN(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6132_ (.A1(_1338_),
    .A2(_2138_),
    .ZN(_2146_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6133_ (.A1(_1653_),
    .A2(_2132_),
    .ZN(_2147_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6134_ (.A1(_1056_),
    .A2(_2146_),
    .A3(_2147_),
    .ZN(_2148_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6135_ (.A1(_1102_),
    .A2(_1513_),
    .B1(_1815_),
    .B2(_3228_),
    .C(_1258_),
    .ZN(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6136_ (.A1(_2066_),
    .A2(_2145_),
    .B1(_2148_),
    .B2(_2149_),
    .ZN(_2150_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6137_ (.I(_1512_),
    .Z(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6138_ (.A1(_1269_),
    .A2(_2110_),
    .ZN(_2152_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6139_ (.A1(_1269_),
    .A2(_2110_),
    .ZN(_2153_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6140_ (.A1(_2112_),
    .A2(_2152_),
    .B(_2153_),
    .ZN(_2154_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6141_ (.A1(_0481_),
    .A2(_0407_),
    .Z(_2155_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6142_ (.A1(_2154_),
    .A2(_2155_),
    .Z(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6143_ (.A1(_2056_),
    .A2(_2156_),
    .ZN(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6144_ (.A1(_1235_),
    .A2(_2151_),
    .B(_2019_),
    .C(_2157_),
    .ZN(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6145_ (.A1(_2000_),
    .A2(_2150_),
    .B(_2158_),
    .ZN(_2159_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6146_ (.A1(_1999_),
    .A2(_2159_),
    .ZN(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6147_ (.A1(\as2650.stack[7][5] ),
    .A2(_1968_),
    .B1(_1975_),
    .B2(\as2650.stack[5][5] ),
    .ZN(_2161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6148_ (.A1(\as2650.stack[6][5] ),
    .A2(_1969_),
    .B1(_2027_),
    .B2(\as2650.stack[4][5] ),
    .ZN(_2162_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6149_ (.A1(_2024_),
    .A2(_2161_),
    .A3(_2162_),
    .ZN(_2163_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6150_ (.I(_1967_),
    .Z(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6151_ (.A1(\as2650.stack[3][5] ),
    .A2(_2164_),
    .B1(_1976_),
    .B2(\as2650.stack[0][5] ),
    .ZN(_2165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6152_ (.A1(\as2650.stack[2][5] ),
    .A2(_1969_),
    .B1(_1975_),
    .B2(\as2650.stack[1][5] ),
    .ZN(_2166_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6153_ (.A1(_2030_),
    .A2(_2165_),
    .A3(_2166_),
    .ZN(_2167_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6154_ (.A1(_2163_),
    .A2(_2167_),
    .ZN(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6155_ (.A1(_1743_),
    .A2(_2132_),
    .B1(_2168_),
    .B2(_1919_),
    .ZN(_2169_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6156_ (.A1(_2139_),
    .A2(_2160_),
    .B(_2169_),
    .ZN(_2170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6157_ (.A1(_2132_),
    .A2(_2140_),
    .B1(_2170_),
    .B2(_2037_),
    .ZN(_2171_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6158_ (.A1(_2130_),
    .A2(_2171_),
    .B(_2039_),
    .ZN(_2172_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6159_ (.A1(_0718_),
    .A2(_1984_),
    .B(_2172_),
    .ZN(_0189_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6160_ (.I(_0720_),
    .Z(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6161_ (.A1(_2141_),
    .A2(_2131_),
    .ZN(_2174_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6162_ (.A1(_2173_),
    .A2(_2174_),
    .Z(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6163_ (.I(_1888_),
    .Z(_2176_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6164_ (.A1(\as2650.pc[6] ),
    .A2(net7),
    .ZN(_2177_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6165_ (.I(_2177_),
    .Z(_2178_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6166_ (.A1(\as2650.pc[4] ),
    .A2(net5),
    .B1(_0481_),
    .B2(_0715_),
    .ZN(_2179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6167_ (.A1(_0716_),
    .A2(_0482_),
    .B(_2179_),
    .ZN(_2180_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6168_ (.A1(_2136_),
    .A2(_2134_),
    .B(_2180_),
    .ZN(_2181_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6169_ (.A1(_2178_),
    .A2(_2181_),
    .ZN(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6170_ (.A1(_2095_),
    .A2(_2175_),
    .B1(_2182_),
    .B2(_2101_),
    .C(_1995_),
    .ZN(_2183_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6171_ (.I(_1799_),
    .Z(_2184_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6172_ (.A1(_2176_),
    .A2(_2183_),
    .B(_2184_),
    .ZN(_2185_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6173_ (.A1(_1099_),
    .A2(_0407_),
    .Z(_2186_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6174_ (.A1(_2154_),
    .A2(_2155_),
    .B(_2186_),
    .ZN(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6175_ (.A1(_0558_),
    .A2(_0486_),
    .Z(_2188_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6176_ (.A1(_2187_),
    .A2(_2188_),
    .B(_2151_),
    .ZN(_2189_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6177_ (.A1(_2187_),
    .A2(_2188_),
    .B(_2189_),
    .ZN(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6178_ (.I(_1562_),
    .Z(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6179_ (.A1(_0559_),
    .A2(_2191_),
    .B(_2020_),
    .ZN(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6180_ (.A1(_2173_),
    .A2(_2142_),
    .Z(_2193_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6181_ (.A1(_2007_),
    .A2(_2182_),
    .ZN(_2194_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6182_ (.A1(_1433_),
    .A2(_2175_),
    .ZN(_2195_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6183_ (.A1(_1890_),
    .A2(_2194_),
    .A3(_2195_),
    .ZN(_2196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6184_ (.A1(_1348_),
    .A2(_1513_),
    .B1(_1815_),
    .B2(_3229_),
    .C(_1210_),
    .ZN(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6185_ (.A1(_2066_),
    .A2(_2193_),
    .B1(_2196_),
    .B2(_2197_),
    .ZN(_2198_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6186_ (.A1(_2190_),
    .A2(_2192_),
    .B1(_2198_),
    .B2(_2065_),
    .ZN(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6187_ (.A1(_1812_),
    .A2(_2199_),
    .ZN(_2200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6188_ (.I(_1742_),
    .Z(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6189_ (.I(_1472_),
    .Z(_2202_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6190_ (.A1(\as2650.stack[7][6] ),
    .A2(_2164_),
    .B1(_1977_),
    .B2(\as2650.stack[6][6] ),
    .ZN(_2203_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6191_ (.A1(\as2650.stack[5][6] ),
    .A2(_1975_),
    .B1(_2079_),
    .B2(\as2650.stack[4][6] ),
    .ZN(_2204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6192_ (.A1(_2203_),
    .A2(_2204_),
    .ZN(_2205_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6193_ (.I(_1967_),
    .Z(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6194_ (.A1(\as2650.stack[3][6] ),
    .A2(_2206_),
    .B1(_0781_),
    .B2(\as2650.stack[1][6] ),
    .ZN(_2207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6195_ (.A1(\as2650.stack[2][6] ),
    .A2(_1924_),
    .B1(_0805_),
    .B2(\as2650.stack[0][6] ),
    .ZN(_2208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6196_ (.I(_1472_),
    .Z(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6197_ (.A1(_2207_),
    .A2(_2208_),
    .B(_2209_),
    .ZN(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6198_ (.I(_1749_),
    .Z(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6199_ (.A1(_2202_),
    .A2(_2205_),
    .B(_2210_),
    .C(_2211_),
    .ZN(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6200_ (.A1(_2201_),
    .A2(_2175_),
    .B(_2212_),
    .ZN(_2213_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6201_ (.A1(_2183_),
    .A2(_2200_),
    .B(_2213_),
    .ZN(_2214_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6202_ (.I(_1800_),
    .Z(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6203_ (.A1(_2175_),
    .A2(_2185_),
    .B1(_2214_),
    .B2(_2215_),
    .ZN(_2216_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6204_ (.I(_1469_),
    .Z(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6205_ (.A1(_2130_),
    .A2(_2216_),
    .B(_2217_),
    .ZN(_2218_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6206_ (.A1(_0722_),
    .A2(_1936_),
    .B(_2218_),
    .ZN(_0190_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6207_ (.I(\as2650.pc[7] ),
    .Z(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6208_ (.I(_1799_),
    .Z(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6209_ (.A1(_0720_),
    .A2(_0715_),
    .A3(_2131_),
    .ZN(_2221_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6210_ (.A1(_0724_),
    .A2(_2221_),
    .Z(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6211_ (.A1(\as2650.pc[7] ),
    .A2(_0557_),
    .ZN(_2223_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6212_ (.A1(_0720_),
    .A2(_0557_),
    .ZN(_2224_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6213_ (.A1(_2178_),
    .A2(_2181_),
    .B(_2224_),
    .ZN(_2225_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6214_ (.A1(_2223_),
    .A2(_2225_),
    .Z(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6215_ (.A1(_1913_),
    .A2(_2226_),
    .ZN(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6216_ (.A1(_1912_),
    .A2(_2222_),
    .B(_2227_),
    .C(_1587_),
    .ZN(_2228_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6217_ (.I(_2228_),
    .ZN(_2229_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6218_ (.I(_1908_),
    .Z(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6219_ (.A1(_0721_),
    .A2(_2142_),
    .ZN(_2231_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6220_ (.A1(_0725_),
    .A2(_2231_),
    .Z(_2232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6221_ (.I(_1126_),
    .Z(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6222_ (.A1(_0659_),
    .A2(_1806_),
    .ZN(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6223_ (.A1(_1268_),
    .A2(_1416_),
    .ZN(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6224_ (.A1(_2233_),
    .A2(_2234_),
    .A3(_2235_),
    .ZN(_2236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6225_ (.A1(_1652_),
    .A2(_2222_),
    .ZN(_2237_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6226_ (.A1(_2009_),
    .A2(_2226_),
    .B(_2237_),
    .C(_3222_),
    .ZN(_2238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6227_ (.A1(_2236_),
    .A2(_2238_),
    .ZN(_2239_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6228_ (.A1(_2230_),
    .A2(_2232_),
    .B1(_2239_),
    .B2(_1310_),
    .ZN(_2240_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6229_ (.A1(_2065_),
    .A2(_2240_),
    .ZN(_2241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6230_ (.A1(_1280_),
    .A2(_0486_),
    .ZN(_2242_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6231_ (.A1(_2187_),
    .A2(_2188_),
    .B(_2242_),
    .ZN(_2243_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6232_ (.A1(net8),
    .A2(_3321_),
    .Z(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6233_ (.A1(_2243_),
    .A2(_2244_),
    .ZN(_2245_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6234_ (.A1(_2243_),
    .A2(_2244_),
    .ZN(_2246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6235_ (.A1(_1807_),
    .A2(_2246_),
    .ZN(_2247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _6236_ (.A1(_1307_),
    .A2(_2013_),
    .B1(_2245_),
    .B2(_2247_),
    .C(_2053_),
    .ZN(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6237_ (.A1(_2064_),
    .A2(_2241_),
    .A3(_2248_),
    .ZN(_2249_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6238_ (.A1(\as2650.stack[5][7] ),
    .A2(_2025_),
    .B1(_2027_),
    .B2(\as2650.stack[4][7] ),
    .C1(\as2650.stack[7][7] ),
    .C2(_0650_),
    .ZN(_2250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6239_ (.A1(\as2650.stack[6][7] ),
    .A2(_1925_),
    .B(_2030_),
    .ZN(_2251_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6240_ (.I(_1970_),
    .Z(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6241_ (.I(_1971_),
    .Z(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6242_ (.A1(\as2650.stack[3][7] ),
    .A2(_0649_),
    .B1(_1924_),
    .B2(\as2650.stack[2][7] ),
    .ZN(_2254_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6243_ (.I(_2254_),
    .ZN(_2255_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6244_ (.A1(\as2650.stack[1][7] ),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[0][7] ),
    .C(_2255_),
    .ZN(_2256_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6245_ (.A1(_2250_),
    .A2(_2251_),
    .B1(_2256_),
    .B2(_1922_),
    .ZN(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6246_ (.A1(_2229_),
    .A2(_2249_),
    .B1(_2257_),
    .B2(_2211_),
    .ZN(_2258_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6247_ (.A1(_1889_),
    .A2(_2229_),
    .B(_1918_),
    .C(_1800_),
    .ZN(_2259_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6248_ (.I(_2222_),
    .ZN(_2260_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6249_ (.A1(_2220_),
    .A2(_2258_),
    .B1(_2259_),
    .B2(_2260_),
    .C(_1886_),
    .ZN(_2261_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6250_ (.A1(_2219_),
    .A2(_1883_),
    .B(_2261_),
    .ZN(_2262_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6251_ (.A1(_1773_),
    .A2(_2262_),
    .ZN(_0191_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6252_ (.A1(_0724_),
    .A2(_2221_),
    .ZN(_2263_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6253_ (.A1(_0729_),
    .A2(_2263_),
    .ZN(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6254_ (.A1(\as2650.pc[8] ),
    .A2(_0558_),
    .Z(_2265_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6255_ (.I(_2265_),
    .ZN(_2266_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6256_ (.A1(_2177_),
    .A2(_2223_),
    .ZN(_2267_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6257_ (.A1(\as2650.pc[7] ),
    .A2(_1211_),
    .B1(_2180_),
    .B2(_2267_),
    .ZN(_2268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6258_ (.A1(_2224_),
    .A2(_2268_),
    .ZN(_2269_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6259_ (.A1(_2134_),
    .A2(_2267_),
    .ZN(_2270_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6260_ (.A1(_2043_),
    .A2(_2096_),
    .A3(_2098_),
    .A4(_2270_),
    .ZN(_2271_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6261_ (.A1(_2269_),
    .A2(_2271_),
    .Z(_2272_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6262_ (.A1(_2266_),
    .A2(_2272_),
    .Z(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6263_ (.A1(_1963_),
    .A2(_2273_),
    .ZN(_2274_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6264_ (.A1(_1940_),
    .A2(_2264_),
    .B(_2274_),
    .C(_1465_),
    .ZN(_2275_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6265_ (.I(\as2650.addr_buff[0] ),
    .ZN(_2276_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6266_ (.A1(_0609_),
    .A2(_3321_),
    .Z(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6267_ (.A1(_2243_),
    .A2(_2244_),
    .B(_2277_),
    .ZN(_2278_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6268_ (.A1(_0687_),
    .A2(_2278_),
    .Z(_2279_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6269_ (.A1(_2276_),
    .A2(_1806_),
    .A3(_2278_),
    .ZN(_2280_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6270_ (.A1(_2276_),
    .A2(_2279_),
    .B(_2280_),
    .ZN(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6271_ (.A1(_2219_),
    .A2(_2231_),
    .ZN(_2282_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6272_ (.A1(_0729_),
    .A2(_2282_),
    .Z(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6273_ (.A1(_1891_),
    .A2(_1453_),
    .ZN(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6274_ (.A1(_1903_),
    .A2(_2284_),
    .ZN(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6275_ (.A1(_1652_),
    .A2(_2273_),
    .ZN(_2286_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6276_ (.A1(_1898_),
    .A2(_2264_),
    .B(_2286_),
    .C(_1145_),
    .ZN(_2287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6277_ (.A1(_1780_),
    .A2(_2285_),
    .B(_2287_),
    .ZN(_2288_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6278_ (.A1(_2230_),
    .A2(_2283_),
    .B1(_2288_),
    .B2(_1075_),
    .ZN(_2289_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6279_ (.A1(_2054_),
    .A2(_2281_),
    .B1(_2289_),
    .B2(_1424_),
    .ZN(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6280_ (.A1(_2064_),
    .A2(_2290_),
    .ZN(_2291_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6281_ (.A1(\as2650.stack[1][8] ),
    .A2(_2082_),
    .B1(_2084_),
    .B2(\as2650.stack[0][8] ),
    .ZN(_2292_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6282_ (.A1(\as2650.stack[3][8] ),
    .A2(_2206_),
    .B1(_2122_),
    .B2(\as2650.stack[2][8] ),
    .ZN(_2293_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6283_ (.A1(_1921_),
    .A2(_2292_),
    .A3(_2293_),
    .ZN(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6284_ (.A1(\as2650.stack[6][8] ),
    .A2(_2122_),
    .B1(_2082_),
    .B2(\as2650.stack[5][8] ),
    .ZN(_2295_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6285_ (.A1(\as2650.stack[7][8] ),
    .A2(_2206_),
    .B1(_2084_),
    .B2(\as2650.stack[4][8] ),
    .ZN(_2296_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6286_ (.A1(_2209_),
    .A2(_2295_),
    .A3(_2296_),
    .ZN(_2297_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6287_ (.A1(_1029_),
    .A2(_2294_),
    .A3(_2297_),
    .ZN(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6288_ (.A1(_1818_),
    .A2(_2264_),
    .B(_2298_),
    .C(_1587_),
    .ZN(_2299_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6289_ (.A1(_2275_),
    .A2(_2291_),
    .B(_2299_),
    .ZN(_2300_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6290_ (.A1(_2176_),
    .A2(_2275_),
    .B(_2184_),
    .ZN(_2301_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6291_ (.A1(_2220_),
    .A2(_2300_),
    .B1(_2301_),
    .B2(_2264_),
    .C(_1886_),
    .ZN(_2302_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6292_ (.A1(_0730_),
    .A2(_1985_),
    .B(_2302_),
    .ZN(_2303_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6293_ (.A1(_1773_),
    .A2(_2303_),
    .ZN(_0192_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6294_ (.I(\as2650.pc[9] ),
    .Z(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6295_ (.A1(_0728_),
    .A2(_2263_),
    .ZN(_2305_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6296_ (.A1(_2304_),
    .A2(_2305_),
    .Z(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6297_ (.A1(_0733_),
    .A2(_1211_),
    .Z(_2307_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6298_ (.I(_2307_),
    .Z(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6299_ (.A1(_0728_),
    .A2(_1280_),
    .ZN(_2309_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6300_ (.A1(_2266_),
    .A2(_2272_),
    .ZN(_2310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6301_ (.A1(_2309_),
    .A2(_2310_),
    .ZN(_2311_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6302_ (.A1(_2308_),
    .A2(_2311_),
    .Z(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6303_ (.A1(_1914_),
    .A2(_2312_),
    .Z(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6304_ (.A1(_1990_),
    .A2(_2306_),
    .B(_2313_),
    .C(_1966_),
    .ZN(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6305_ (.A1(_2176_),
    .A2(_2314_),
    .B(_2184_),
    .ZN(_2315_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6306_ (.A1(_1540_),
    .A2(_2280_),
    .Z(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6307_ (.A1(_0728_),
    .A2(_2219_),
    .A3(_2231_),
    .ZN(_2317_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6308_ (.A1(_2304_),
    .A2(_2317_),
    .Z(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6309_ (.A1(_2007_),
    .A2(_2312_),
    .ZN(_2319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6310_ (.A1(_2009_),
    .A2(_2306_),
    .B(_2233_),
    .ZN(_2320_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6311_ (.I(\as2650.addr_buff[1] ),
    .Z(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6312_ (.A1(_2321_),
    .A2(_1453_),
    .ZN(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6313_ (.A1(_1959_),
    .A2(_2322_),
    .ZN(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6314_ (.A1(_2319_),
    .A2(_2320_),
    .B1(_2323_),
    .B2(_1780_),
    .ZN(_2324_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6315_ (.A1(_2066_),
    .A2(_2318_),
    .B1(_2324_),
    .B2(_1310_),
    .ZN(_2325_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6316_ (.A1(_2054_),
    .A2(_2316_),
    .B1(_2325_),
    .B2(_1802_),
    .ZN(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6317_ (.A1(_1812_),
    .A2(_2326_),
    .ZN(_2327_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6318_ (.A1(\as2650.stack[7][9] ),
    .A2(_2164_),
    .B1(_2078_),
    .B2(\as2650.stack[6][9] ),
    .ZN(_2328_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6319_ (.A1(\as2650.stack[5][9] ),
    .A2(_2076_),
    .B1(_2079_),
    .B2(\as2650.stack[4][9] ),
    .ZN(_2329_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6320_ (.A1(_2328_),
    .A2(_2329_),
    .ZN(_2330_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6321_ (.A1(\as2650.stack[2][9] ),
    .A2(_2122_),
    .B1(_0805_),
    .B2(\as2650.stack[0][9] ),
    .ZN(_2331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6322_ (.A1(\as2650.stack[3][9] ),
    .A2(_0649_),
    .B1(_0781_),
    .B2(\as2650.stack[1][9] ),
    .ZN(_2332_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6323_ (.A1(_2331_),
    .A2(_2332_),
    .B(_2209_),
    .ZN(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6324_ (.A1(_2202_),
    .A2(_2330_),
    .B(_2333_),
    .C(_2211_),
    .ZN(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6325_ (.A1(_2201_),
    .A2(_2306_),
    .B(_2334_),
    .ZN(_2335_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6326_ (.A1(_2314_),
    .A2(_2327_),
    .B(_2335_),
    .ZN(_2336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6327_ (.A1(_2306_),
    .A2(_2315_),
    .B1(_2336_),
    .B2(_2215_),
    .ZN(_2337_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6328_ (.A1(_2130_),
    .A2(_2337_),
    .B(_2217_),
    .ZN(_2338_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6329_ (.A1(_0735_),
    .A2(_1936_),
    .B(_2338_),
    .ZN(_0193_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6330_ (.I(\as2650.pc[10] ),
    .Z(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6331_ (.A1(\as2650.pc[9] ),
    .A2(\as2650.pc[8] ),
    .A3(_2263_),
    .ZN(_2340_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6332_ (.A1(_2339_),
    .A2(_2340_),
    .Z(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6333_ (.I(_1211_),
    .Z(_2342_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6334_ (.A1(_0739_),
    .A2(_2342_),
    .Z(_2343_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6335_ (.A1(\as2650.pc[9] ),
    .A2(\as2650.pc[8] ),
    .B(_2342_),
    .ZN(_2344_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6336_ (.A1(_2310_),
    .A2(_2307_),
    .B(_2344_),
    .ZN(_2345_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6337_ (.A1(_2343_),
    .A2(_2345_),
    .Z(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_2 _6338_ (.A1(_2095_),
    .A2(_2341_),
    .B1(_2346_),
    .B2(_2101_),
    .C(_1465_),
    .ZN(_2347_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6339_ (.A1(_2176_),
    .A2(_2347_),
    .B(_2184_),
    .ZN(_2348_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6340_ (.I(_2321_),
    .ZN(_2349_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6341_ (.A1(_2276_),
    .A2(_2349_),
    .A3(_1744_),
    .A4(_2278_),
    .ZN(_2350_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6342_ (.A1(_1542_),
    .A2(_2350_),
    .Z(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6343_ (.A1(_0734_),
    .A2(_2317_),
    .ZN(_2352_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6344_ (.A1(_0740_),
    .A2(_2352_),
    .Z(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6345_ (.A1(_2003_),
    .A2(_0687_),
    .B(_2018_),
    .ZN(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6346_ (.A1(_1780_),
    .A2(_2354_),
    .B(_1210_),
    .ZN(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6347_ (.A1(_2007_),
    .A2(_2346_),
    .ZN(_2356_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6348_ (.A1(_1433_),
    .A2(_2341_),
    .ZN(_2357_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6349_ (.A1(_1890_),
    .A2(_2356_),
    .A3(_2357_),
    .ZN(_2358_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6350_ (.A1(_2230_),
    .A2(_2353_),
    .B1(_2355_),
    .B2(_2358_),
    .ZN(_2359_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6351_ (.A1(_2054_),
    .A2(_2351_),
    .B1(_2359_),
    .B2(_1802_),
    .ZN(_2360_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6352_ (.A1(_1812_),
    .A2(_2360_),
    .ZN(_2361_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6353_ (.A1(\as2650.stack[6][10] ),
    .A2(_1977_),
    .B1(_1976_),
    .B2(\as2650.stack[4][10] ),
    .ZN(_2362_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6354_ (.A1(\as2650.stack[7][10] ),
    .A2(_2164_),
    .B1(_2076_),
    .B2(\as2650.stack[5][10] ),
    .ZN(_2363_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6355_ (.A1(_2362_),
    .A2(_2363_),
    .ZN(_2364_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6356_ (.A1(\as2650.stack[3][10] ),
    .A2(_2206_),
    .B1(_0781_),
    .B2(\as2650.stack[1][10] ),
    .ZN(_2365_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6357_ (.A1(\as2650.stack[2][10] ),
    .A2(_1924_),
    .B1(_0805_),
    .B2(\as2650.stack[0][10] ),
    .ZN(_2366_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6358_ (.A1(_2365_),
    .A2(_2366_),
    .B(_2209_),
    .ZN(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6359_ (.A1(_2202_),
    .A2(_2364_),
    .B(_2367_),
    .C(_1749_),
    .ZN(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6360_ (.A1(_2201_),
    .A2(_2341_),
    .B(_2368_),
    .ZN(_2369_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6361_ (.A1(_2347_),
    .A2(_2361_),
    .B(_2369_),
    .ZN(_2370_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6362_ (.A1(_2341_),
    .A2(_2348_),
    .B1(_2370_),
    .B2(_2215_),
    .ZN(_2371_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6363_ (.A1(_2130_),
    .A2(_2371_),
    .B(_2217_),
    .ZN(_2372_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6364_ (.A1(_0741_),
    .A2(_1936_),
    .B(_2372_),
    .ZN(_0194_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6365_ (.I(_2339_),
    .Z(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6366_ (.A1(_2373_),
    .A2(_2352_),
    .ZN(_2374_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6367_ (.A1(_0744_),
    .A2(_2374_),
    .Z(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6368_ (.A1(_0739_),
    .A2(_2340_),
    .ZN(_2376_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6369_ (.A1(\as2650.pc[11] ),
    .A2(_2376_),
    .Z(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6370_ (.I(_2377_),
    .Z(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6371_ (.A1(_1909_),
    .A2(_2375_),
    .B1(_2378_),
    .B2(_1775_),
    .ZN(_2379_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6372_ (.A1(_0743_),
    .A2(_2342_),
    .Z(_2380_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6373_ (.A1(_2339_),
    .A2(_1212_),
    .ZN(_2381_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6374_ (.A1(_2339_),
    .A2(_2342_),
    .Z(_2382_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6375_ (.A1(_2382_),
    .A2(_2345_),
    .ZN(_2383_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6376_ (.A1(_2381_),
    .A2(_2383_),
    .ZN(_2384_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6377_ (.A1(_2380_),
    .A2(_2384_),
    .ZN(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6378_ (.A1(_1652_),
    .A2(_2377_),
    .Z(_2386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6379_ (.A1(_1338_),
    .A2(_2385_),
    .B(_2386_),
    .C(_2233_),
    .ZN(_2387_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6380_ (.A1(_1298_),
    .A2(_1562_),
    .B(_2233_),
    .ZN(_2388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6381_ (.A1(\as2650.addr_buff[3] ),
    .A2(_1512_),
    .B(_2388_),
    .ZN(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6382_ (.A1(_1566_),
    .A2(_1424_),
    .A3(_2387_),
    .A4(_2389_),
    .Z(_2390_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6383_ (.A1(_1802_),
    .A2(_2379_),
    .B(_2390_),
    .ZN(_2391_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _6384_ (.I(\as2650.addr_buff[3] ),
    .ZN(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_2 _6385_ (.A1(\as2650.addr_buff[0] ),
    .A2(_2321_),
    .A3(\as2650.addr_buff[2] ),
    .ZN(_2393_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6386_ (.A1(_0686_),
    .A2(_2278_),
    .A3(_2393_),
    .ZN(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6387_ (.A1(_2392_),
    .A2(_2394_),
    .Z(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6388_ (.A1(_1781_),
    .A2(_2377_),
    .ZN(_2396_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6389_ (.A1(_1781_),
    .A2(_2395_),
    .B(_2396_),
    .C(_1639_),
    .ZN(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6390_ (.A1(_1999_),
    .A2(_2391_),
    .A3(_2397_),
    .ZN(_2398_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6391_ (.A1(_1990_),
    .A2(_2378_),
    .B1(_2385_),
    .B2(_1915_),
    .C(_1463_),
    .ZN(_2399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6392_ (.A1(\as2650.stack[5][11] ),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[4][11] ),
    .ZN(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6393_ (.A1(\as2650.stack[7][11] ),
    .A2(_0650_),
    .B1(_0754_),
    .B2(\as2650.stack[6][11] ),
    .ZN(_2401_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6394_ (.A1(_1473_),
    .A2(_2400_),
    .A3(_2401_),
    .ZN(_2402_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _6395_ (.A1(\as2650.stack[1][11] ),
    .A2(_2025_),
    .B1(_2027_),
    .B2(\as2650.stack[0][11] ),
    .C1(\as2650.stack[2][11] ),
    .C2(_0754_),
    .ZN(_2403_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6396_ (.A1(\as2650.stack[3][11] ),
    .A2(_1929_),
    .B(_2202_),
    .ZN(_2404_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6397_ (.A1(_2403_),
    .A2(_2404_),
    .B(_2211_),
    .ZN(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6398_ (.A1(_2201_),
    .A2(_2378_),
    .B1(_2402_),
    .B2(_2405_),
    .ZN(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6399_ (.A1(_2398_),
    .A2(_2399_),
    .B(_2406_),
    .ZN(_2407_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6400_ (.A1(_1801_),
    .A2(_2407_),
    .ZN(_2408_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6401_ (.A1(_1885_),
    .A2(_2378_),
    .B(_1935_),
    .ZN(_2409_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6402_ (.A1(_0744_),
    .A2(_1883_),
    .B1(_2408_),
    .B2(_2409_),
    .C(_1853_),
    .ZN(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6403_ (.A1(_1545_),
    .A2(_2394_),
    .Z(_2410_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6404_ (.A1(_1542_),
    .A2(_1545_),
    .A3(_1548_),
    .A4(_2350_),
    .ZN(_2411_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6405_ (.A1(_1548_),
    .A2(_2410_),
    .B(_2411_),
    .C(_2020_),
    .ZN(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6406_ (.I(\as2650.pc[11] ),
    .Z(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6407_ (.A1(_2413_),
    .A2(_2376_),
    .ZN(_2414_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6408_ (.A1(_0747_),
    .A2(_2414_),
    .Z(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6409_ (.I(_2415_),
    .ZN(_2416_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6410_ (.A1(_2413_),
    .A2(_2373_),
    .A3(_2352_),
    .ZN(_2417_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6411_ (.A1(_0747_),
    .A2(_2417_),
    .Z(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6412_ (.A1(_1649_),
    .A2(_2230_),
    .A3(_2418_),
    .ZN(_2419_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6413_ (.A1(_2310_),
    .A2(_2308_),
    .ZN(_2420_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6414_ (.A1(_2343_),
    .A2(_2380_),
    .ZN(_2421_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6415_ (.A1(_0743_),
    .A2(_0558_),
    .B(_2381_),
    .C(_2344_),
    .ZN(_2422_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6416_ (.A1(_2420_),
    .A2(_2421_),
    .B(_2422_),
    .ZN(_2423_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6417_ (.A1(\as2650.pc[12] ),
    .A2(_1280_),
    .Z(_2424_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6418_ (.A1(_2423_),
    .A2(_2424_),
    .Z(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6419_ (.A1(_1898_),
    .A2(_2415_),
    .ZN(_2426_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6420_ (.A1(_1653_),
    .A2(_2425_),
    .B(_2426_),
    .C(_1435_),
    .ZN(_2427_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6421_ (.A1(\as2650.addr_buff[4] ),
    .A2(_2004_),
    .ZN(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6422_ (.A1(_1134_),
    .A2(_2114_),
    .A3(_2428_),
    .ZN(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6423_ (.A1(_1310_),
    .A2(_1431_),
    .A3(_2427_),
    .A4(_2429_),
    .ZN(_2430_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6424_ (.A1(_1889_),
    .A2(_2416_),
    .B(_2419_),
    .C(_2430_),
    .ZN(_2431_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6425_ (.A1(_1914_),
    .A2(_2425_),
    .ZN(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6426_ (.A1(_1912_),
    .A2(_2415_),
    .B1(_2431_),
    .B2(_1776_),
    .C(_2432_),
    .ZN(_2433_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6427_ (.A1(_2412_),
    .A2(_2433_),
    .B(_2088_),
    .ZN(_2434_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6428_ (.A1(\as2650.stack[5][12] ),
    .A2(_2252_),
    .B1(_2253_),
    .B2(\as2650.stack[4][12] ),
    .ZN(_2435_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6429_ (.A1(\as2650.stack[7][12] ),
    .A2(_1929_),
    .B1(_0754_),
    .B2(\as2650.stack[6][12] ),
    .ZN(_2436_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6430_ (.A1(_1473_),
    .A2(_2435_),
    .A3(_2436_),
    .ZN(_2437_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6431_ (.A1(\as2650.stack[3][12] ),
    .A2(_1929_),
    .B1(_2252_),
    .B2(\as2650.stack[1][12] ),
    .ZN(_2438_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6432_ (.A1(\as2650.stack[2][12] ),
    .A2(_1925_),
    .B1(_2253_),
    .B2(\as2650.stack[0][12] ),
    .ZN(_2439_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6433_ (.A1(_1922_),
    .A2(_2438_),
    .A3(_2439_),
    .ZN(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6434_ (.A1(_1919_),
    .A2(_2437_),
    .A3(_2440_),
    .ZN(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6435_ (.A1(_1918_),
    .A2(_2416_),
    .B(_2441_),
    .ZN(_2442_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6436_ (.A1(_2434_),
    .A2(_2442_),
    .B(_1801_),
    .ZN(_2443_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6437_ (.A1(_1885_),
    .A2(_2415_),
    .B(_1935_),
    .ZN(_2444_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6438_ (.A1(_0748_),
    .A2(_1883_),
    .B1(_2443_),
    .B2(_2444_),
    .C(_1595_),
    .ZN(_0196_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6439_ (.I(_1744_),
    .Z(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6440_ (.I(_2445_),
    .Z(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6441_ (.I(_2446_),
    .Z(_2447_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6442_ (.I(_1500_),
    .Z(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6443_ (.I(_2448_),
    .Z(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6444_ (.I(_2449_),
    .Z(_2450_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6445_ (.A1(_2450_),
    .A2(_3391_),
    .ZN(_2451_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6446_ (.I(_1685_),
    .Z(_2452_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6447_ (.A1(_2452_),
    .A2(_3302_),
    .ZN(_2453_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6448_ (.A1(_2447_),
    .A2(_2451_),
    .A3(_2453_),
    .ZN(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6449_ (.I(_1125_),
    .Z(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6450_ (.A1(_2056_),
    .A2(_3431_),
    .B(_2455_),
    .ZN(_2456_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6451_ (.I(_1263_),
    .Z(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6452_ (.I(_1218_),
    .Z(_2458_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6453_ (.I(_1091_),
    .Z(_2459_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6454_ (.A1(\as2650.psu[0] ),
    .A2(_2459_),
    .ZN(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6455_ (.I(_1873_),
    .Z(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6456_ (.A1(\as2650.carry ),
    .A2(_2461_),
    .B(_2458_),
    .ZN(_2462_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6457_ (.A1(_2458_),
    .A2(_3343_),
    .B1(_2460_),
    .B2(_2462_),
    .ZN(_2463_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6458_ (.A1(_1225_),
    .A2(_2463_),
    .ZN(_2464_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6459_ (.I(_1088_),
    .Z(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6460_ (.A1(_2465_),
    .A2(_0892_),
    .B(_1264_),
    .ZN(_2466_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6461_ (.A1(_1488_),
    .A2(_2457_),
    .B1(_2464_),
    .B2(_2466_),
    .ZN(_2467_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _6462_ (.A1(_3433_),
    .A2(_1426_),
    .A3(_1597_),
    .B(_1678_),
    .ZN(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6463_ (.A1(_1124_),
    .A2(_3285_),
    .ZN(_2469_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6464_ (.A1(_3256_),
    .A2(_1530_),
    .B(_2469_),
    .ZN(_2470_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6465_ (.A1(_1183_),
    .A2(_0920_),
    .B1(_1618_),
    .B2(_1420_),
    .C(_2470_),
    .ZN(_2471_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6466_ (.A1(_1132_),
    .A2(_3314_),
    .A3(_3230_),
    .ZN(_2472_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6467_ (.A1(_0673_),
    .A2(_1558_),
    .A3(_1176_),
    .A4(_2472_),
    .Z(_2473_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6468_ (.A1(_3265_),
    .A2(_0920_),
    .B(_1152_),
    .C(_1158_),
    .ZN(_2474_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6469_ (.A1(_2471_),
    .A2(_2473_),
    .A3(_2474_),
    .ZN(_2475_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6470_ (.I(_3306_),
    .Z(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6471_ (.A1(_3184_),
    .A2(_2476_),
    .A3(_1129_),
    .ZN(_2477_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6472_ (.A1(_3303_),
    .A2(_0379_),
    .A3(_1168_),
    .A4(_1657_),
    .ZN(_2478_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_2 _6473_ (.A1(_1052_),
    .A2(_1065_),
    .A3(_1086_),
    .A4(_1121_),
    .ZN(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6474_ (.A1(_3174_),
    .A2(_3316_),
    .A3(_3262_),
    .ZN(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6475_ (.A1(_1506_),
    .A2(_1342_),
    .A3(_2480_),
    .ZN(_2481_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6476_ (.I(_1502_),
    .Z(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6477_ (.A1(_1123_),
    .A2(_2482_),
    .B1(_1520_),
    .B2(_0658_),
    .ZN(_2483_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6478_ (.A1(_2481_),
    .A2(_2483_),
    .ZN(_2484_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6479_ (.A1(_1138_),
    .A2(_2478_),
    .B(_2479_),
    .C(_2484_),
    .ZN(_2485_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6480_ (.A1(_0896_),
    .A2(_0881_),
    .A3(_1151_),
    .ZN(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6481_ (.A1(_0913_),
    .A2(_3188_),
    .A3(_3382_),
    .A4(_0916_),
    .ZN(_2487_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6482_ (.A1(_2486_),
    .A2(_2487_),
    .B(_0869_),
    .ZN(_2488_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _6483_ (.A1(_1172_),
    .A2(_2477_),
    .A3(_2485_),
    .A4(_2488_),
    .ZN(_2489_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6484_ (.A1(_2468_),
    .A2(_2475_),
    .A3(_2489_),
    .ZN(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6485_ (.I(_2490_),
    .Z(_2491_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6486_ (.A1(_3370_),
    .A2(_1524_),
    .B1(_1850_),
    .B2(_3548_),
    .C(_2491_),
    .ZN(_2492_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6487_ (.A1(_2454_),
    .A2(_2456_),
    .B1(_2467_),
    .B2(_1583_),
    .C(_2492_),
    .ZN(_2493_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6488_ (.I(_2490_),
    .Z(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6489_ (.A1(_3311_),
    .A2(_2494_),
    .B(_1736_),
    .ZN(_2495_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6490_ (.A1(_2493_),
    .A2(_2495_),
    .ZN(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6491_ (.I(_1115_),
    .Z(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6492_ (.I(_2490_),
    .Z(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6493_ (.A1(_3483_),
    .A2(_2497_),
    .ZN(_2498_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6494_ (.I(_2445_),
    .Z(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6495_ (.A1(_1685_),
    .A2(_3492_),
    .ZN(_2500_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6496_ (.A1(_1764_),
    .A2(_3449_),
    .ZN(_2501_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6497_ (.A1(_2499_),
    .A2(_2500_),
    .A3(_2501_),
    .ZN(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6498_ (.A1(_2056_),
    .A2(_3524_),
    .B(_2455_),
    .ZN(_2503_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6499_ (.A1(_1966_),
    .A2(_3476_),
    .ZN(_2504_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6500_ (.I(_1091_),
    .Z(_2505_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6501_ (.A1(_1279_),
    .A2(_1091_),
    .ZN(_2506_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6502_ (.A1(\as2650.psu[1] ),
    .A2(_2505_),
    .B(_2506_),
    .C(_1090_),
    .ZN(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6503_ (.A1(_3283_),
    .A2(_3451_),
    .B1(_0332_),
    .B2(_1088_),
    .C(_1263_),
    .ZN(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6504_ (.A1(_1292_),
    .A2(_1232_),
    .B1(_2507_),
    .B2(_2508_),
    .C(_1587_),
    .ZN(_2509_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6505_ (.A1(_1834_),
    .A2(_2504_),
    .A3(_2509_),
    .ZN(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6506_ (.A1(_2491_),
    .A2(_2510_),
    .ZN(_2511_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6507_ (.A1(_0892_),
    .A2(_1855_),
    .B1(_2502_),
    .B2(_2503_),
    .C(_2511_),
    .ZN(_2512_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6508_ (.A1(_2496_),
    .A2(_2498_),
    .A3(_2512_),
    .ZN(_0198_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6509_ (.A1(_0438_),
    .A2(_3582_),
    .ZN(_2513_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6510_ (.A1(_0268_),
    .A2(_0272_),
    .ZN(_2514_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6511_ (.A1(_2513_),
    .A2(_2514_),
    .ZN(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6512_ (.I(_1201_),
    .Z(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6513_ (.I(_1763_),
    .Z(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6514_ (.A1(_2449_),
    .A2(_3571_),
    .ZN(_2518_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6515_ (.A1(_2517_),
    .A2(_3577_),
    .B(_2518_),
    .C(_2446_),
    .ZN(_2519_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6516_ (.A1(_2499_),
    .A2(_2515_),
    .B(_2516_),
    .C(_2519_),
    .ZN(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6517_ (.A1(\as2650.psu[2] ),
    .A2(_2505_),
    .Z(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6518_ (.A1(\as2650.overflow ),
    .A2(_2461_),
    .B(_2521_),
    .C(_1312_),
    .ZN(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6519_ (.A1(_2458_),
    .A2(_3529_),
    .B1(_0976_),
    .B2(_1225_),
    .C(_2522_),
    .ZN(_2523_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6520_ (.A1(_3543_),
    .A2(_1229_),
    .B(_1078_),
    .ZN(_2524_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6521_ (.A1(_1229_),
    .A2(_2523_),
    .B(_2524_),
    .ZN(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6522_ (.A1(_3556_),
    .A2(_1779_),
    .B1(_1854_),
    .B2(_0332_),
    .ZN(_2526_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6523_ (.A1(_2497_),
    .A2(_2520_),
    .A3(_2525_),
    .A4(_2526_),
    .Z(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6524_ (.A1(_1710_),
    .A2(_2494_),
    .B(_1736_),
    .ZN(_2528_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6525_ (.A1(_2527_),
    .A2(_2528_),
    .ZN(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6526_ (.A1(_2517_),
    .A2(_0331_),
    .ZN(_2529_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6527_ (.A1(_1685_),
    .A2(_0325_),
    .ZN(_2530_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6528_ (.A1(_2499_),
    .A2(_2529_),
    .A3(_2530_),
    .ZN(_2531_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6529_ (.A1(_2447_),
    .A2(_0315_),
    .B(_2516_),
    .C(_2531_),
    .ZN(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6530_ (.I(\as2650.psu[3] ),
    .ZN(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6531_ (.A1(_2533_),
    .A2(_2505_),
    .B(_1090_),
    .ZN(_2534_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6532_ (.A1(_3319_),
    .A2(_1092_),
    .B(_2534_),
    .ZN(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6533_ (.A1(_2458_),
    .A2(_0332_),
    .B1(_0477_),
    .B2(_1225_),
    .C(_3212_),
    .ZN(_2536_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6534_ (.A1(_1544_),
    .A2(_1229_),
    .B1(_2535_),
    .B2(_2536_),
    .C(_1078_),
    .ZN(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6535_ (.A1(_1628_),
    .A2(_1779_),
    .B1(_1854_),
    .B2(_3537_),
    .C(_2537_),
    .ZN(_2538_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _6536_ (.A1(_2497_),
    .A2(_2532_),
    .A3(_2538_),
    .Z(_2539_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6537_ (.A1(_0354_),
    .A2(_2494_),
    .B(_1461_),
    .ZN(_2540_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6538_ (.A1(_2539_),
    .A2(_2540_),
    .ZN(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6539_ (.I(_2446_),
    .Z(_2541_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6540_ (.I(_1201_),
    .Z(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6541_ (.A1(_2450_),
    .A2(_0406_),
    .ZN(_2543_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6542_ (.A1(_2452_),
    .A2(_0400_),
    .ZN(_2544_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6543_ (.A1(_2541_),
    .A2(_2543_),
    .A3(_2544_),
    .ZN(_2545_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6544_ (.A1(_2541_),
    .A2(_0394_),
    .B(_2542_),
    .C(_2545_),
    .ZN(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6545_ (.A1(_0422_),
    .A2(_1837_),
    .ZN(_2547_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6546_ (.A1(_0477_),
    .A2(_1854_),
    .ZN(_2548_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6547_ (.A1(_1288_),
    .A2(_2461_),
    .ZN(_2549_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6548_ (.A1(_3432_),
    .A2(_2461_),
    .B(_2549_),
    .C(_1312_),
    .ZN(_2550_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6549_ (.A1(_1220_),
    .A2(_3537_),
    .B1(_0549_),
    .B2(_1223_),
    .ZN(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6550_ (.A1(_2550_),
    .A2(_2551_),
    .B(_1264_),
    .ZN(_2552_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6551_ (.A1(_1720_),
    .A2(_2457_),
    .B(_1583_),
    .C(_2552_),
    .ZN(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6552_ (.A1(_2497_),
    .A2(_2547_),
    .A3(_2548_),
    .A4(_2553_),
    .Z(_2554_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6553_ (.I(_2490_),
    .Z(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6554_ (.A1(_0975_),
    .A2(_2555_),
    .B(_2217_),
    .ZN(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6555_ (.A1(_2546_),
    .A2(_2554_),
    .B(_2556_),
    .ZN(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6556_ (.A1(_1519_),
    .A2(_0505_),
    .Z(_2557_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6557_ (.A1(_1764_),
    .A2(_0475_),
    .B(_2557_),
    .C(_2499_),
    .ZN(_2558_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6558_ (.A1(_2013_),
    .A2(_0466_),
    .B(_2516_),
    .C(_2558_),
    .ZN(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6559_ (.A1(_1466_),
    .A2(_0480_),
    .ZN(_2560_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6560_ (.I(_1049_),
    .Z(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6561_ (.A1(\as2650.psl[5] ),
    .A2(_2459_),
    .B(_2561_),
    .ZN(_2562_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6562_ (.A1(_1296_),
    .A2(_1092_),
    .B(_2562_),
    .ZN(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6563_ (.A1(_1218_),
    .A2(_0477_),
    .ZN(_2564_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6564_ (.A1(_2465_),
    .A2(_0604_),
    .B(_2564_),
    .C(_1232_),
    .ZN(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6565_ (.A1(_1103_),
    .A2(_2457_),
    .B1(_2563_),
    .B2(_2565_),
    .C(_2088_),
    .ZN(_2566_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6566_ (.A1(_1741_),
    .A2(_2560_),
    .A3(_2566_),
    .ZN(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6567_ (.A1(_0549_),
    .A2(_1850_),
    .B(_2559_),
    .C(_2567_),
    .ZN(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6568_ (.I(_1469_),
    .Z(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6569_ (.A1(_0476_),
    .A2(_2555_),
    .B(_2569_),
    .ZN(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6570_ (.A1(_2494_),
    .A2(_2568_),
    .B(_2570_),
    .ZN(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6571_ (.A1(_2450_),
    .A2(_0546_),
    .ZN(_2571_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6572_ (.A1(_2452_),
    .A2(_0569_),
    .ZN(_2572_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6573_ (.A1(_2447_),
    .A2(_2571_),
    .A3(_2572_),
    .ZN(_2573_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6574_ (.A1(_2541_),
    .A2(_0537_),
    .B(_2542_),
    .C(_2573_),
    .ZN(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6575_ (.A1(_1117_),
    .A2(_2505_),
    .B(_2561_),
    .ZN(_2575_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6576_ (.A1(net24),
    .A2(_2459_),
    .B(_2575_),
    .ZN(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6577_ (.I(_0574_),
    .Z(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6578_ (.A1(_1223_),
    .A2(_2577_),
    .B1(_0549_),
    .B2(_1220_),
    .ZN(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6579_ (.A1(_2576_),
    .A2(_2578_),
    .B(_1232_),
    .ZN(_2579_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6580_ (.A1(_1349_),
    .A2(_2457_),
    .B(_1583_),
    .C(_2579_),
    .ZN(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6581_ (.A1(_2491_),
    .A2(_2580_),
    .ZN(_2581_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6582_ (.A1(_0556_),
    .A2(_1837_),
    .B1(_1855_),
    .B2(_0989_),
    .C(_2581_),
    .ZN(_2582_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6583_ (.A1(_1728_),
    .A2(_2555_),
    .B(_2569_),
    .ZN(_2583_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6584_ (.A1(_2574_),
    .A2(_2582_),
    .B(_2583_),
    .ZN(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6585_ (.A1(_2450_),
    .A2(_0603_),
    .ZN(_2584_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6586_ (.A1(_2452_),
    .A2(_0623_),
    .ZN(_2585_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6587_ (.A1(_2447_),
    .A2(_2584_),
    .A3(_2585_),
    .ZN(_2586_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6588_ (.A1(_2541_),
    .A2(_0597_),
    .B(_2542_),
    .C(_2586_),
    .ZN(_2587_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6589_ (.A1(_1254_),
    .A2(_2459_),
    .B(_2561_),
    .ZN(_2588_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6590_ (.A1(_1295_),
    .A2(_1092_),
    .B(_2588_),
    .ZN(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6591_ (.A1(_1351_),
    .A2(_1264_),
    .B1(_1265_),
    .B2(_2589_),
    .C(_1516_),
    .ZN(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6592_ (.A1(_2491_),
    .A2(_2590_),
    .ZN(_2591_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6593_ (.A1(_0607_),
    .A2(_1837_),
    .B1(_1855_),
    .B2(_2577_),
    .C(_2591_),
    .ZN(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6594_ (.A1(_0617_),
    .A2(_2555_),
    .B(_2569_),
    .ZN(_2593_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6595_ (.A1(_2587_),
    .A2(_2592_),
    .B(_2593_),
    .ZN(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6596_ (.A1(_0689_),
    .A2(_0755_),
    .ZN(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6597_ (.I(_2594_),
    .Z(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6598_ (.I(_2595_),
    .Z(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6599_ (.I(_2594_),
    .Z(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6600_ (.A1(\as2650.stack[7][0] ),
    .A2(_2597_),
    .ZN(_2598_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6601_ (.A1(_0835_),
    .A2(_2596_),
    .B(_2598_),
    .ZN(_0205_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6602_ (.A1(\as2650.stack[7][1] ),
    .A2(_2597_),
    .ZN(_2599_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6603_ (.A1(_0841_),
    .A2(_2596_),
    .B(_2599_),
    .ZN(_0206_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6604_ (.A1(\as2650.stack[7][2] ),
    .A2(_2597_),
    .ZN(_2600_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6605_ (.A1(_0701_),
    .A2(_2596_),
    .B(_2600_),
    .ZN(_0207_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6606_ (.A1(\as2650.stack[7][3] ),
    .A2(_2597_),
    .ZN(_2601_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6607_ (.A1(_0705_),
    .A2(_2596_),
    .B(_2601_),
    .ZN(_0208_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6608_ (.I(_2595_),
    .Z(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6609_ (.I(_2594_),
    .Z(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6610_ (.A1(\as2650.stack[7][4] ),
    .A2(_2603_),
    .ZN(_2604_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6611_ (.A1(_0710_),
    .A2(_2602_),
    .B(_2604_),
    .ZN(_0209_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6612_ (.A1(\as2650.stack[7][5] ),
    .A2(_2603_),
    .ZN(_2605_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6613_ (.A1(_0717_),
    .A2(_2602_),
    .B(_2605_),
    .ZN(_0210_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6614_ (.A1(\as2650.stack[7][6] ),
    .A2(_2603_),
    .ZN(_2606_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6615_ (.A1(_0721_),
    .A2(_2602_),
    .B(_2606_),
    .ZN(_0211_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6616_ (.A1(\as2650.stack[7][7] ),
    .A2(_2603_),
    .ZN(_2607_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6617_ (.A1(_0850_),
    .A2(_2602_),
    .B(_2607_),
    .ZN(_0212_));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _6618_ (.I0(_0852_),
    .I1(\as2650.stack[7][8] ),
    .S(_2595_),
    .Z(_2608_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6619_ (.I(_2608_),
    .Z(_0213_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6620_ (.I(_2595_),
    .Z(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6621_ (.I(_2594_),
    .Z(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6622_ (.A1(\as2650.stack[7][9] ),
    .A2(_2610_),
    .ZN(_2611_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6623_ (.A1(_0734_),
    .A2(_2609_),
    .B(_2611_),
    .ZN(_0214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6624_ (.A1(\as2650.stack[7][10] ),
    .A2(_2610_),
    .ZN(_2612_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6625_ (.A1(_0740_),
    .A2(_2609_),
    .B(_2612_),
    .ZN(_0215_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6626_ (.A1(\as2650.stack[7][11] ),
    .A2(_2610_),
    .ZN(_2613_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6627_ (.A1(_0858_),
    .A2(_2609_),
    .B(_2613_),
    .ZN(_0216_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6628_ (.A1(\as2650.stack[7][12] ),
    .A2(_2610_),
    .ZN(_2614_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6629_ (.A1(_0860_),
    .A2(_2609_),
    .B(_2614_),
    .ZN(_0217_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6630_ (.A1(_1508_),
    .A2(_1510_),
    .ZN(_2615_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6631_ (.A1(_1558_),
    .A2(_2615_),
    .ZN(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6632_ (.A1(_0665_),
    .A2(_1506_),
    .A3(_1612_),
    .ZN(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6633_ (.A1(_2616_),
    .A2(_2617_),
    .B(_1067_),
    .C(_1326_),
    .ZN(_2618_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _6634_ (.A1(_1526_),
    .A2(_1869_),
    .A3(_1604_),
    .A4(_1874_),
    .ZN(_2619_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _6635_ (.A1(_1615_),
    .A2(_1670_),
    .A3(_1868_),
    .A4(_2619_),
    .Z(_2620_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6636_ (.A1(_1602_),
    .A2(_2620_),
    .ZN(_2621_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6637_ (.A1(_1632_),
    .A2(_2618_),
    .A3(_2621_),
    .ZN(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6638_ (.I(_2622_),
    .Z(_2623_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6639_ (.I(_2623_),
    .Z(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6640_ (.I(_2624_),
    .Z(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6641_ (.I(_1498_),
    .Z(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6642_ (.I(_1503_),
    .Z(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6643_ (.I(_2627_),
    .Z(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6644_ (.I(_3187_),
    .Z(_2629_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6645_ (.A1(_2629_),
    .A2(_3302_),
    .ZN(_2630_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6646_ (.A1(_0879_),
    .A2(_2630_),
    .Z(_2631_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6647_ (.A1(_0658_),
    .A2(_3230_),
    .ZN(_2632_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6648_ (.I(_2632_),
    .Z(_2633_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6649_ (.A1(_3391_),
    .A2(_2633_),
    .ZN(_2634_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6650_ (.A1(_0879_),
    .A2(_2634_),
    .Z(_2635_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6651_ (.A1(_2628_),
    .A2(_2631_),
    .B1(_2635_),
    .B2(_2517_),
    .ZN(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6652_ (.I(net25),
    .Z(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6653_ (.I(_1617_),
    .Z(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6654_ (.I(_2638_),
    .Z(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6655_ (.I(_1125_),
    .Z(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6656_ (.A1(_2637_),
    .A2(_2639_),
    .B1(_1828_),
    .B2(_1896_),
    .C(_2640_),
    .ZN(_2641_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6657_ (.A1(_2626_),
    .A2(_2636_),
    .B(_2641_),
    .ZN(_2642_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6658_ (.A1(_1455_),
    .A2(_3236_),
    .ZN(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6659_ (.I(_2643_),
    .Z(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6660_ (.A1(_1134_),
    .A2(_1511_),
    .ZN(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6661_ (.A1(_2637_),
    .A2(_1807_),
    .B(_1894_),
    .ZN(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6662_ (.A1(_1344_),
    .A2(_1896_),
    .B1(_2645_),
    .B2(_2646_),
    .ZN(_2647_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6663_ (.A1(_1146_),
    .A2(_1811_),
    .B(_2643_),
    .ZN(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6664_ (.A1(_2644_),
    .A2(_2647_),
    .B1(_2648_),
    .B2(_0645_),
    .ZN(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6665_ (.A1(_1785_),
    .A2(_2649_),
    .ZN(_2650_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6666_ (.A1(_2642_),
    .A2(_2650_),
    .ZN(_2651_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6667_ (.A1(_1850_),
    .A2(_1689_),
    .ZN(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6668_ (.A1(_1634_),
    .A2(_2651_),
    .B1(_2652_),
    .B2(_1897_),
    .ZN(_2653_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6669_ (.I(_2623_),
    .Z(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6670_ (.A1(_2637_),
    .A2(_2654_),
    .B(_2569_),
    .ZN(_2655_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6671_ (.A1(_2625_),
    .A2(_2653_),
    .B(_2655_),
    .ZN(_0218_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6672_ (.I(_1589_),
    .Z(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6673_ (.A1(_1162_),
    .A2(_2656_),
    .ZN(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6674_ (.I(_2657_),
    .Z(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6675_ (.I(_1501_),
    .Z(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6676_ (.A1(net52),
    .A2(_2637_),
    .Z(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6677_ (.A1(_1527_),
    .A2(_2626_),
    .ZN(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6678_ (.I(_2476_),
    .Z(_2662_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6679_ (.A1(_3372_),
    .A2(_3301_),
    .ZN(_2663_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6680_ (.A1(_3465_),
    .A2(_3492_),
    .A3(_2663_),
    .Z(_2664_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6681_ (.I(_3307_),
    .Z(_2665_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6682_ (.A1(_1238_),
    .A2(_2665_),
    .ZN(_2666_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6683_ (.I(_2627_),
    .Z(_2667_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6684_ (.A1(_2662_),
    .A2(_2664_),
    .B(_2666_),
    .C(_2667_),
    .ZN(_2668_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6685_ (.A1(\as2650.addr_buff[7] ),
    .A2(_3230_),
    .Z(_2669_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6686_ (.I(_2669_),
    .Z(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6687_ (.I(_2670_),
    .Z(_2671_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6688_ (.A1(_3372_),
    .A2(_3390_),
    .ZN(_2672_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6689_ (.A1(_3465_),
    .A2(_3449_),
    .A3(_2672_),
    .Z(_2673_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6690_ (.I(_2669_),
    .Z(_2674_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6691_ (.A1(_1238_),
    .A2(_2674_),
    .ZN(_2675_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6692_ (.A1(_2671_),
    .A2(_2673_),
    .B(_2675_),
    .C(_2448_),
    .ZN(_2676_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6693_ (.A1(_2668_),
    .A2(_2676_),
    .ZN(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6694_ (.A1(_2661_),
    .A2(_2677_),
    .ZN(_2678_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6695_ (.A1(_2659_),
    .A2(_2660_),
    .B(_2678_),
    .C(_1787_),
    .ZN(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6696_ (.I(_1831_),
    .Z(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6697_ (.A1(_0642_),
    .A2(net1),
    .ZN(_2681_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6698_ (.A1(_2681_),
    .A2(_1947_),
    .Z(_2682_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6699_ (.A1(_2680_),
    .A2(_2682_),
    .B(_2640_),
    .ZN(_2683_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6700_ (.I(_2648_),
    .Z(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6701_ (.A1(_3222_),
    .A2(_1811_),
    .ZN(_2685_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6702_ (.A1(_1807_),
    .A2(_2660_),
    .ZN(_2686_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6703_ (.A1(_1944_),
    .A2(_2686_),
    .ZN(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6704_ (.A1(_1327_),
    .A2(_1948_),
    .B1(_2685_),
    .B2(_2687_),
    .ZN(_2688_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6705_ (.I(_2688_),
    .ZN(_2689_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6706_ (.A1(_1937_),
    .A2(_2684_),
    .B1(_2689_),
    .B2(_2644_),
    .ZN(_2690_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6707_ (.A1(_2679_),
    .A2(_2683_),
    .B1(_2690_),
    .B2(_1205_),
    .ZN(_2691_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6708_ (.I(_2656_),
    .Z(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6709_ (.A1(_1937_),
    .A2(_2658_),
    .B1(_2691_),
    .B2(_2692_),
    .ZN(_2693_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6710_ (.I(_1459_),
    .Z(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6711_ (.A1(net52),
    .A2(_2654_),
    .B(_2694_),
    .ZN(_2695_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6712_ (.A1(_2625_),
    .A2(_2693_),
    .B(_2695_),
    .ZN(_0219_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6713_ (.I(_2623_),
    .Z(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6714_ (.A1(net52),
    .A2(net25),
    .ZN(_2697_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6715_ (.A1(net27),
    .A2(_2697_),
    .Z(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6716_ (.A1(_2681_),
    .A2(_1947_),
    .B(_1992_),
    .ZN(_2699_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6717_ (.A1(_1991_),
    .A2(_2699_),
    .Z(_2700_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6718_ (.I(_1676_),
    .Z(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6719_ (.A1(_3462_),
    .A2(_3491_),
    .ZN(_2702_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6720_ (.A1(_3463_),
    .A2(_3491_),
    .ZN(_2703_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6721_ (.A1(_2663_),
    .A2(_2702_),
    .B(_2703_),
    .ZN(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6722_ (.A1(_1239_),
    .A2(_3577_),
    .Z(_2705_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6723_ (.A1(_2704_),
    .A2(_2705_),
    .B(_3307_),
    .ZN(_2706_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6724_ (.A1(_2704_),
    .A2(_2705_),
    .B(_2706_),
    .ZN(_2707_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6725_ (.A1(_1241_),
    .A2(_2629_),
    .B(_2627_),
    .C(_2707_),
    .ZN(_2708_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6726_ (.A1(_3463_),
    .A2(_3448_),
    .ZN(_2709_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6727_ (.A1(_3463_),
    .A2(_3448_),
    .ZN(_2710_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6728_ (.A1(_2672_),
    .A2(_2709_),
    .B(_2710_),
    .ZN(_2711_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6729_ (.A1(_3541_),
    .A2(_3571_),
    .Z(_2712_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6730_ (.A1(_2711_),
    .A2(_2712_),
    .B(_2670_),
    .ZN(_2713_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6731_ (.A1(_2711_),
    .A2(_2712_),
    .B(_2713_),
    .ZN(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6732_ (.I(_1500_),
    .Z(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6733_ (.A1(_1240_),
    .A2(_2632_),
    .B(_2714_),
    .C(_2715_),
    .ZN(_2716_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6734_ (.A1(_2708_),
    .A2(_2716_),
    .ZN(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6735_ (.A1(_2701_),
    .A2(_2717_),
    .ZN(_2718_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6736_ (.A1(_1501_),
    .A2(_2698_),
    .B1(_2700_),
    .B2(_1786_),
    .C(_2718_),
    .ZN(_2719_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6737_ (.A1(_1434_),
    .A2(_0357_),
    .ZN(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6738_ (.A1(_1056_),
    .A2(_1344_),
    .B(_2720_),
    .ZN(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6739_ (.A1(_2004_),
    .A2(_2698_),
    .B(_2005_),
    .ZN(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6740_ (.A1(_2065_),
    .A2(_2010_),
    .B1(_2685_),
    .B2(_2722_),
    .ZN(_2723_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6741_ (.A1(_0700_),
    .A2(_2721_),
    .B1(_2723_),
    .B2(_2720_),
    .ZN(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6742_ (.A1(_1201_),
    .A2(_2719_),
    .B1(_2724_),
    .B2(_1834_),
    .ZN(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6743_ (.I(_2622_),
    .Z(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6744_ (.A1(_0701_),
    .A2(_2657_),
    .B1(_2725_),
    .B2(_2656_),
    .C(_2726_),
    .ZN(_2727_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6745_ (.A1(net27),
    .A2(_2696_),
    .B(_2727_),
    .ZN(_2728_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6746_ (.A1(_1772_),
    .A2(_2728_),
    .ZN(_0220_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6747_ (.A1(_2046_),
    .A2(_2699_),
    .ZN(_2729_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6748_ (.A1(_0700_),
    .A2(_3543_),
    .B(_2729_),
    .ZN(_2730_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6749_ (.A1(_2045_),
    .A2(_2730_),
    .Z(_2731_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6750_ (.A1(net27),
    .A2(net26),
    .A3(net25),
    .ZN(_2732_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6751_ (.A1(net28),
    .A2(_2732_),
    .Z(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6752_ (.A1(_3573_),
    .A2(_3576_),
    .B(_3540_),
    .ZN(_2734_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6753_ (.A1(_3540_),
    .A2(_3573_),
    .A3(_3576_),
    .ZN(_2735_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6754_ (.A1(_2704_),
    .A2(_2734_),
    .B(_2735_),
    .ZN(_2736_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6755_ (.A1(_0344_),
    .A2(_0325_),
    .A3(_2736_),
    .Z(_2737_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6756_ (.A1(_0345_),
    .A2(_2476_),
    .ZN(_2738_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6757_ (.A1(_2665_),
    .A2(_2737_),
    .B(_2738_),
    .C(_2667_),
    .ZN(_2739_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6758_ (.A1(_1298_),
    .A2(_0331_),
    .Z(_2740_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _6759_ (.A1(_3566_),
    .A2(_3570_),
    .B(_3541_),
    .ZN(_2741_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_2 _6760_ (.A1(_3540_),
    .A2(_3566_),
    .A3(_3570_),
    .ZN(_2742_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6761_ (.A1(_2711_),
    .A2(_2741_),
    .B(_2742_),
    .ZN(_2743_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6762_ (.A1(_2740_),
    .A2(_2743_),
    .B(_2670_),
    .ZN(_2744_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6763_ (.A1(_2740_),
    .A2(_2743_),
    .B(_2744_),
    .ZN(_2745_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6764_ (.A1(_1544_),
    .A2(_2633_),
    .B(_2745_),
    .C(_2448_),
    .ZN(_2746_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6765_ (.I(_1677_),
    .Z(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6766_ (.A1(_2739_),
    .A2(_2746_),
    .B(_2747_),
    .ZN(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6767_ (.A1(_2638_),
    .A2(_2733_),
    .B(_2748_),
    .C(_1828_),
    .ZN(_2749_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6768_ (.A1(_2680_),
    .A2(_2731_),
    .B(_2749_),
    .ZN(_2750_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6769_ (.A1(_1242_),
    .A2(_2191_),
    .ZN(_2751_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6770_ (.A1(_1418_),
    .A2(_2733_),
    .B(_2751_),
    .ZN(_2752_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6771_ (.A1(_2041_),
    .A2(_2684_),
    .B1(_2752_),
    .B2(_1428_),
    .C(_1257_),
    .ZN(_2753_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6772_ (.A1(_2542_),
    .A2(_2750_),
    .B1(_2753_),
    .B2(_2050_),
    .ZN(_2754_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6773_ (.A1(_2041_),
    .A2(_2658_),
    .B1(_2754_),
    .B2(_2692_),
    .ZN(_2755_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6774_ (.A1(net28),
    .A2(_2654_),
    .B(_2694_),
    .ZN(_2756_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6775_ (.A1(_2625_),
    .A2(_2755_),
    .B(_2756_),
    .ZN(_0221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6776_ (.A1(_2046_),
    .A2(_2699_),
    .B(_2044_),
    .C(_2047_),
    .ZN(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6777_ (.A1(_2043_),
    .A2(_2757_),
    .ZN(_2758_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6778_ (.A1(_2097_),
    .A2(_2758_),
    .Z(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6779_ (.I(net28),
    .ZN(_2760_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6780_ (.A1(_2760_),
    .A2(_2732_),
    .ZN(_2761_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6781_ (.A1(net29),
    .A2(_2761_),
    .Z(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _6782_ (.I(_0343_),
    .Z(_2763_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6783_ (.A1(_2763_),
    .A2(_0324_),
    .ZN(_2764_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6784_ (.A1(_2763_),
    .A2(_0324_),
    .B1(_2704_),
    .B2(_2734_),
    .C(_2735_),
    .ZN(_2765_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6785_ (.A1(_2764_),
    .A2(_2765_),
    .ZN(_2766_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6786_ (.A1(_0424_),
    .A2(_0400_),
    .A3(_2766_),
    .Z(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6787_ (.A1(_2629_),
    .A2(_2767_),
    .ZN(_2768_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6788_ (.A1(_1719_),
    .A2(_2629_),
    .B(_2667_),
    .C(_2768_),
    .ZN(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6789_ (.A1(_2763_),
    .A2(_0330_),
    .ZN(_2770_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6790_ (.A1(_1270_),
    .A2(_0406_),
    .Z(_2771_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_4 _6791_ (.A1(_2763_),
    .A2(_0330_),
    .B1(_2711_),
    .B2(_2741_),
    .C(_2742_),
    .ZN(_2772_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6792_ (.A1(_2770_),
    .A2(_2771_),
    .A3(_2772_),
    .ZN(_2773_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6793_ (.A1(_2770_),
    .A2(_2772_),
    .B(_2771_),
    .ZN(_2774_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6794_ (.A1(_2633_),
    .A2(_2774_),
    .ZN(_2775_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6795_ (.A1(_1719_),
    .A2(_2633_),
    .B1(_2773_),
    .B2(_2775_),
    .C(_1763_),
    .ZN(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6796_ (.A1(_2769_),
    .A2(_2776_),
    .B(_2626_),
    .ZN(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6797_ (.A1(_1832_),
    .A2(_2759_),
    .B1(_2762_),
    .B2(_2639_),
    .C(_2777_),
    .ZN(_2778_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6798_ (.A1(_1417_),
    .A2(_2762_),
    .ZN(_2779_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6799_ (.A1(_1234_),
    .A2(_1429_),
    .B(_2779_),
    .ZN(_2780_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6800_ (.A1(_2645_),
    .A2(_2780_),
    .ZN(_2781_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6801_ (.A1(_2064_),
    .A2(_2100_),
    .B(_2781_),
    .ZN(_2782_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6802_ (.A1(_2135_),
    .A2(_2721_),
    .B1(_2782_),
    .B2(_2720_),
    .C(_1204_),
    .ZN(_2783_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6803_ (.A1(_2455_),
    .A2(_2778_),
    .B(_2783_),
    .ZN(_2784_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6804_ (.A1(_2135_),
    .A2(_2652_),
    .B1(_2784_),
    .B2(_1634_),
    .ZN(_2785_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6805_ (.I(_2623_),
    .Z(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6806_ (.A1(net29),
    .A2(_2786_),
    .B(_2694_),
    .ZN(_2787_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6807_ (.A1(_2625_),
    .A2(_2785_),
    .B(_2787_),
    .ZN(_0222_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6808_ (.I(_2657_),
    .Z(_2788_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6809_ (.A1(_2097_),
    .A2(_2758_),
    .ZN(_2789_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6810_ (.A1(_0710_),
    .A2(_0425_),
    .B(_2789_),
    .ZN(_2790_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6811_ (.A1(_2134_),
    .A2(_2790_),
    .Z(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6812_ (.A1(net29),
    .A2(_2761_),
    .Z(_2792_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6813_ (.A1(net51),
    .A2(_2792_),
    .ZN(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6814_ (.A1(_1269_),
    .A2(_0399_),
    .ZN(_2794_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6815_ (.A1(_0423_),
    .A2(_0399_),
    .ZN(_2795_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6816_ (.A1(_2764_),
    .A2(_2794_),
    .A3(_2765_),
    .B(_2795_),
    .ZN(_2796_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6817_ (.A1(_0483_),
    .A2(_0475_),
    .A3(_2796_),
    .Z(_2797_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6818_ (.A1(_1101_),
    .A2(_2476_),
    .ZN(_2798_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6819_ (.A1(_2665_),
    .A2(_2797_),
    .B(_2798_),
    .C(_2627_),
    .ZN(_2799_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6820_ (.A1(_0423_),
    .A2(_0405_),
    .ZN(_2800_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6821_ (.A1(_0423_),
    .A2(_0405_),
    .ZN(_2801_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_2 _6822_ (.A1(_2770_),
    .A2(_2800_),
    .A3(_2772_),
    .B(_2801_),
    .ZN(_2802_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6823_ (.A1(_0482_),
    .A2(_0505_),
    .A3(_2802_),
    .Z(_2803_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6824_ (.A1(_1101_),
    .A2(_2674_),
    .ZN(_2804_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6825_ (.A1(_2674_),
    .A2(_2803_),
    .B(_2804_),
    .C(_2715_),
    .ZN(_2805_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6826_ (.A1(_2799_),
    .A2(_2805_),
    .B(_1677_),
    .ZN(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6827_ (.A1(_2638_),
    .A2(_2793_),
    .B(_2806_),
    .C(_1831_),
    .ZN(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6828_ (.A1(_2680_),
    .A2(_2791_),
    .B(_2807_),
    .C(_2640_),
    .ZN(_2808_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6829_ (.A1(_1689_),
    .A2(_2808_),
    .ZN(_2809_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6830_ (.A1(_1102_),
    .A2(_2191_),
    .ZN(_2810_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6831_ (.A1(_1418_),
    .A2(_2793_),
    .B(_2810_),
    .ZN(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6832_ (.A1(_2141_),
    .A2(_2648_),
    .B1(_2811_),
    .B2(_1428_),
    .ZN(_2812_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6833_ (.A1(_1915_),
    .A2(_2138_),
    .B(_2812_),
    .C(_2220_),
    .ZN(_2813_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6834_ (.A1(_2141_),
    .A2(_2788_),
    .B(_2809_),
    .C(_2813_),
    .ZN(_2814_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6835_ (.A1(net51),
    .A2(_2726_),
    .ZN(_2815_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6836_ (.A1(_2696_),
    .A2(_2814_),
    .B(_2815_),
    .C(_1691_),
    .ZN(_0223_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6837_ (.I(_2726_),
    .Z(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6838_ (.A1(_2133_),
    .A2(_2789_),
    .ZN(_2817_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6839_ (.A1(_2180_),
    .A2(_2817_),
    .ZN(_2818_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6840_ (.A1(_2178_),
    .A2(_2818_),
    .Z(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6841_ (.A1(net51),
    .A2(_2792_),
    .ZN(_2820_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6842_ (.A1(net32),
    .A2(_2820_),
    .Z(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6843_ (.A1(_1099_),
    .A2(_0474_),
    .Z(_2822_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6844_ (.A1(_1099_),
    .A2(_0474_),
    .Z(_2823_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_4 _6845_ (.A1(_2796_),
    .A2(_2822_),
    .B(_2823_),
    .ZN(_2824_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6846_ (.A1(_1272_),
    .A2(_0568_),
    .A3(_2824_),
    .Z(_2825_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6847_ (.A1(_1348_),
    .A2(_2665_),
    .ZN(_2826_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6848_ (.A1(_2662_),
    .A2(_2825_),
    .B(_2826_),
    .C(_2667_),
    .ZN(_2827_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6849_ (.A1(_1100_),
    .A2(_0504_),
    .Z(_2828_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6850_ (.A1(_1100_),
    .A2(_0504_),
    .Z(_2829_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6851_ (.A1(_2828_),
    .A2(_2802_),
    .B(_2829_),
    .ZN(_2830_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6852_ (.A1(_1272_),
    .A2(_0545_),
    .A3(_2830_),
    .Z(_2831_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6853_ (.A1(_1348_),
    .A2(_2674_),
    .ZN(_2832_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6854_ (.A1(_2671_),
    .A2(_2831_),
    .B(_2832_),
    .C(_2448_),
    .ZN(_2833_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6855_ (.A1(_2827_),
    .A2(_2833_),
    .B(_2747_),
    .ZN(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6856_ (.A1(_2638_),
    .A2(_2821_),
    .B(_2834_),
    .C(_1828_),
    .ZN(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6857_ (.A1(_1832_),
    .A2(_2819_),
    .B(_2835_),
    .C(_2455_),
    .ZN(_2836_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6858_ (.I(_2648_),
    .Z(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6859_ (.A1(_1429_),
    .A2(_2821_),
    .ZN(_2838_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6860_ (.A1(_1349_),
    .A2(_1418_),
    .B(_2838_),
    .ZN(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6861_ (.A1(_1776_),
    .A2(_2182_),
    .B1(_2645_),
    .B2(_2839_),
    .ZN(_2840_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6862_ (.A1(_2173_),
    .A2(_2837_),
    .B1(_2840_),
    .B2(_2644_),
    .C(_1257_),
    .ZN(_2841_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6863_ (.A1(_2836_),
    .A2(_2841_),
    .B(_1689_),
    .ZN(_2842_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6864_ (.A1(_2173_),
    .A2(_2658_),
    .B(_2842_),
    .ZN(_2843_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6865_ (.A1(net32),
    .A2(_2786_),
    .B(_2694_),
    .ZN(_2844_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6866_ (.A1(_2816_),
    .A2(_2843_),
    .B(_2844_),
    .ZN(_0224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6867_ (.A1(_1213_),
    .A2(_0568_),
    .ZN(_2845_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6868_ (.A1(_1213_),
    .A2(_0569_),
    .ZN(_2846_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6869_ (.A1(_2845_),
    .A2(_2824_),
    .B(_2846_),
    .ZN(_2847_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6870_ (.A1(_1553_),
    .A2(_0623_),
    .A3(_2847_),
    .Z(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6871_ (.A1(_1231_),
    .A2(_2662_),
    .ZN(_2849_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6872_ (.A1(_2662_),
    .A2(_2848_),
    .B(_2849_),
    .C(_2628_),
    .ZN(_2850_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6873_ (.A1(_1213_),
    .A2(_0545_),
    .ZN(_2851_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6874_ (.A1(_1272_),
    .A2(_0546_),
    .ZN(_2852_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6875_ (.A1(_2851_),
    .A2(_2830_),
    .B(_2852_),
    .ZN(_2853_));
 gf180mcu_fd_sc_mcu7t5v0__xor3_1 _6876_ (.A1(_1553_),
    .A2(_0603_),
    .A3(_2853_),
    .Z(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6877_ (.A1(_1231_),
    .A2(_2671_),
    .ZN(_2855_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6878_ (.A1(_2671_),
    .A2(_2854_),
    .B(_2855_),
    .C(_2517_),
    .ZN(_2856_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6879_ (.A1(_2850_),
    .A2(_2856_),
    .ZN(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6880_ (.I(net33),
    .ZN(_2858_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6881_ (.A1(net32),
    .A2(net51),
    .A3(_2792_),
    .ZN(_2859_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6882_ (.A1(_2858_),
    .A2(_2859_),
    .Z(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6883_ (.I(_1786_),
    .Z(_2861_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6884_ (.A1(_2659_),
    .A2(_2860_),
    .B(_2861_),
    .ZN(_2862_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6885_ (.A1(_2701_),
    .A2(_2857_),
    .B(_2862_),
    .ZN(_2863_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6886_ (.A1(_2178_),
    .A2(_2818_),
    .B(_2224_),
    .ZN(_2864_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6887_ (.A1(_2223_),
    .A2(_2864_),
    .Z(_2865_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _6888_ (.I(_1683_),
    .Z(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6889_ (.A1(_2861_),
    .A2(_2865_),
    .B(_2866_),
    .ZN(_2867_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6890_ (.A1(_1745_),
    .A2(_2860_),
    .ZN(_2868_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6891_ (.A1(_2235_),
    .A2(_2868_),
    .ZN(_2869_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6892_ (.I(_1428_),
    .Z(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6893_ (.A1(_2219_),
    .A2(_2837_),
    .B1(_2869_),
    .B2(_2870_),
    .C(_2227_),
    .ZN(_2871_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6894_ (.A1(_0725_),
    .A2(_2652_),
    .B1(_2871_),
    .B2(_2215_),
    .ZN(_2872_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6895_ (.A1(_2863_),
    .A2(_2867_),
    .B(_2872_),
    .ZN(_2873_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _6896_ (.I(_1459_),
    .Z(_2874_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6897_ (.A1(net33),
    .A2(_2786_),
    .B(_2874_),
    .ZN(_2875_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6898_ (.A1(_2816_),
    .A2(_2873_),
    .B(_2875_),
    .ZN(_0225_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6899_ (.A1(_2858_),
    .A2(_2859_),
    .ZN(_2876_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6900_ (.A1(net50),
    .A2(_2876_),
    .Z(_2877_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6901_ (.A1(_0610_),
    .A2(_0602_),
    .ZN(_2878_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _6902_ (.A1(_2851_),
    .A2(_2830_),
    .B(_2878_),
    .C(_2852_),
    .ZN(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6903_ (.A1(_1268_),
    .A2(_0602_),
    .ZN(_2880_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6904_ (.A1(_2670_),
    .A2(_2880_),
    .ZN(_2881_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6905_ (.A1(_2879_),
    .A2(_2881_),
    .ZN(_2882_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6906_ (.A1(_1537_),
    .A2(_2882_),
    .Z(_2883_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6907_ (.A1(_0609_),
    .A2(_0622_),
    .ZN(_2884_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_4 _6908_ (.A1(_2845_),
    .A2(_2824_),
    .B(_2884_),
    .C(_2846_),
    .ZN(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6909_ (.A1(_0610_),
    .A2(_0622_),
    .ZN(_2886_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _6910_ (.A1(_3307_),
    .A2(_2886_),
    .ZN(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6911_ (.A1(_2885_),
    .A2(_2887_),
    .ZN(_2888_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6912_ (.A1(_1537_),
    .A2(_2888_),
    .Z(_2889_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6913_ (.A1(_2449_),
    .A2(_2883_),
    .B1(_2889_),
    .B2(_2628_),
    .ZN(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6914_ (.A1(_2659_),
    .A2(_2877_),
    .B1(_2890_),
    .B2(_2747_),
    .ZN(_2891_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6915_ (.A1(_2267_),
    .A2(_2817_),
    .B(_2269_),
    .ZN(_2892_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6916_ (.A1(_2265_),
    .A2(_2892_),
    .ZN(_2893_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6917_ (.A1(_2265_),
    .A2(_2892_),
    .ZN(_2894_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6918_ (.I(_2894_),
    .ZN(_2895_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6919_ (.A1(_2680_),
    .A2(_2893_),
    .A3(_2895_),
    .ZN(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6920_ (.A1(_1847_),
    .A2(_2891_),
    .B(_2896_),
    .C(_2516_),
    .ZN(_2897_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6921_ (.A1(_2445_),
    .A2(_2877_),
    .ZN(_2898_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _6922_ (.A1(_2284_),
    .A2(_2685_),
    .Z(_2899_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6923_ (.A1(_2000_),
    .A2(_2286_),
    .B1(_2898_),
    .B2(_2899_),
    .ZN(_2900_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6924_ (.A1(_0729_),
    .A2(_2721_),
    .B1(_2900_),
    .B2(_2720_),
    .ZN(_2901_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6925_ (.A1(_2220_),
    .A2(_2901_),
    .ZN(_2902_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6926_ (.A1(_0730_),
    .A2(_2788_),
    .B1(_2897_),
    .B2(_2692_),
    .C(_2902_),
    .ZN(_2903_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6927_ (.A1(net50),
    .A2(_2786_),
    .B(_2874_),
    .ZN(_2904_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6928_ (.A1(_2816_),
    .A2(_2903_),
    .B(_2904_),
    .ZN(_0226_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6929_ (.A1(net50),
    .A2(_2876_),
    .ZN(_2905_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6930_ (.A1(net35),
    .A2(_2905_),
    .Z(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6931_ (.A1(_1891_),
    .A2(_2885_),
    .A3(_2887_),
    .ZN(_2907_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6932_ (.A1(_1540_),
    .A2(_2907_),
    .Z(_2908_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6933_ (.A1(_1891_),
    .A2(_2879_),
    .A3(_2881_),
    .ZN(_2909_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6934_ (.A1(_2321_),
    .A2(_2909_),
    .Z(_2910_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6935_ (.A1(_2628_),
    .A2(_2908_),
    .B1(_2910_),
    .B2(_2449_),
    .ZN(_2911_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6936_ (.A1(_2747_),
    .A2(_2911_),
    .ZN(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _6937_ (.A1(_2639_),
    .A2(_2906_),
    .B(_2912_),
    .C(_1847_),
    .ZN(_2913_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6938_ (.A1(_2309_),
    .A2(_2895_),
    .ZN(_2914_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6939_ (.A1(_2308_),
    .A2(_2914_),
    .Z(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6940_ (.A1(_2861_),
    .A2(_2915_),
    .B(_2866_),
    .ZN(_2916_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6941_ (.A1(_2151_),
    .A2(_2906_),
    .B(_2322_),
    .ZN(_2917_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6942_ (.A1(_2304_),
    .A2(_2837_),
    .B1(_2917_),
    .B2(_2870_),
    .C(_1939_),
    .ZN(_2918_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6943_ (.A1(_2313_),
    .A2(_2918_),
    .ZN(_2919_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6944_ (.A1(_2304_),
    .A2(_2788_),
    .B1(_2913_),
    .B2(_2916_),
    .C(_2919_),
    .ZN(_2920_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6945_ (.A1(net35),
    .A2(_2624_),
    .B(_2874_),
    .ZN(_2921_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6946_ (.A1(_2816_),
    .A2(_2920_),
    .B(_2921_),
    .ZN(_0227_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_2 _6947_ (.A1(_2879_),
    .A2(_2881_),
    .B(_1519_),
    .ZN(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6948_ (.A1(_2885_),
    .A2(_2887_),
    .B(_2715_),
    .C(_2482_),
    .ZN(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6949_ (.A1(_1537_),
    .A2(_1540_),
    .B(_2482_),
    .ZN(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__or3_1 _6950_ (.A1(_2922_),
    .A2(_2923_),
    .A3(_2924_),
    .Z(_2925_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6951_ (.A1(_2885_),
    .A2(_2887_),
    .B(_2715_),
    .ZN(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _6952_ (.A1(_2482_),
    .A2(_2393_),
    .Z(_2927_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6953_ (.A1(_2926_),
    .A2(_2922_),
    .A3(_2927_),
    .ZN(_2928_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6954_ (.A1(_2003_),
    .A2(_2925_),
    .B(_2928_),
    .ZN(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _6955_ (.A1(net35),
    .A2(net50),
    .A3(_2876_),
    .ZN(_2930_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6956_ (.A1(net36),
    .A2(_2930_),
    .Z(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6957_ (.A1(_2639_),
    .A2(_2931_),
    .ZN(_2932_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _6958_ (.A1(_2626_),
    .A2(_2929_),
    .B(_2932_),
    .C(_1787_),
    .ZN(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6959_ (.I(_2344_),
    .ZN(_2934_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6960_ (.A1(_2308_),
    .A2(_2895_),
    .ZN(_2935_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6961_ (.A1(_2934_),
    .A2(_2935_),
    .B(_2382_),
    .ZN(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _6962_ (.A1(_2382_),
    .A2(_2934_),
    .A3(_2935_),
    .ZN(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6963_ (.A1(_1786_),
    .A2(_2937_),
    .ZN(_2938_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6964_ (.A1(_2936_),
    .A2(_2938_),
    .B(_2640_),
    .ZN(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6965_ (.A1(_2151_),
    .A2(_2931_),
    .ZN(_2940_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6966_ (.A1(_1542_),
    .A2(_2191_),
    .B(_2940_),
    .ZN(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6967_ (.A1(_1344_),
    .A2(_2346_),
    .B1(_2645_),
    .B2(_2941_),
    .ZN(_2942_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6968_ (.A1(_2373_),
    .A2(_2684_),
    .B1(_2942_),
    .B2(_2644_),
    .ZN(_2943_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6969_ (.A1(_2933_),
    .A2(_2939_),
    .B1(_2943_),
    .B2(_1205_),
    .ZN(_2944_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _6970_ (.A1(_2373_),
    .A2(_2658_),
    .B1(_2944_),
    .B2(_2692_),
    .ZN(_2945_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6971_ (.A1(net36),
    .A2(_2624_),
    .B(_2874_),
    .ZN(_2946_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6972_ (.A1(_2696_),
    .A2(_2945_),
    .B(_2946_),
    .ZN(_0228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6973_ (.A1(_3141_),
    .A2(_1617_),
    .ZN(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_2 _6974_ (.A1(_2947_),
    .A2(_2393_),
    .B(_2922_),
    .C(_2923_),
    .ZN(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _6975_ (.A1(_2392_),
    .A2(_2926_),
    .A3(_2922_),
    .A4(_2927_),
    .Z(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6976_ (.A1(_1545_),
    .A2(_2948_),
    .B(_2949_),
    .ZN(_2950_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _6977_ (.I(net36),
    .ZN(_2951_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6978_ (.A1(_2951_),
    .A2(_2930_),
    .ZN(_2952_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6979_ (.A1(net37),
    .A2(_2952_),
    .Z(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6980_ (.A1(_2659_),
    .A2(_2953_),
    .B(_1787_),
    .ZN(_2954_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6981_ (.A1(_2701_),
    .A2(_2950_),
    .B(_2954_),
    .ZN(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6982_ (.A1(_2381_),
    .A2(_2936_),
    .ZN(_2956_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _6983_ (.A1(_2380_),
    .A2(_2956_),
    .Z(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6984_ (.A1(_2861_),
    .A2(_2957_),
    .B(_2866_),
    .ZN(_2958_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6985_ (.A1(_1963_),
    .A2(_2385_),
    .ZN(_2959_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6986_ (.A1(_2445_),
    .A2(_2953_),
    .ZN(_2960_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6987_ (.A1(_2392_),
    .A2(_2446_),
    .B(_2960_),
    .ZN(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _6988_ (.A1(_2413_),
    .A2(_2837_),
    .B1(_2961_),
    .B2(_2870_),
    .C(_1939_),
    .ZN(_2962_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6989_ (.A1(_2959_),
    .A2(_2962_),
    .ZN(_2963_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _6990_ (.A1(_2413_),
    .A2(_2788_),
    .B1(_2955_),
    .B2(_2958_),
    .C(_2963_),
    .ZN(_2964_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6991_ (.A1(net37),
    .A2(_2624_),
    .B(_1460_),
    .ZN(_2965_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6992_ (.A1(_2696_),
    .A2(_2964_),
    .B(_2965_),
    .ZN(_0229_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _6993_ (.A1(net37),
    .A2(_2952_),
    .ZN(_2966_));
 gf180mcu_fd_sc_mcu7t5v0__xnor2_1 _6994_ (.A1(net38),
    .A2(_2966_),
    .ZN(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _6995_ (.A1(_2947_),
    .A2(_2967_),
    .ZN(_2968_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6996_ (.A1(_2392_),
    .A2(_2947_),
    .B(\as2650.addr_buff[4] ),
    .ZN(_2969_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _6997_ (.A1(_1548_),
    .A2(_2949_),
    .B1(_2948_),
    .B2(_2969_),
    .ZN(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _6998_ (.A1(_2968_),
    .A2(_2970_),
    .B(_2701_),
    .ZN(_2971_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _6999_ (.A1(_2421_),
    .A2(_2935_),
    .B(_2422_),
    .ZN(_2972_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7000_ (.A1(_2424_),
    .A2(_2972_),
    .Z(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7001_ (.A1(_2661_),
    .A2(_2967_),
    .B(_2866_),
    .ZN(_2974_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7002_ (.A1(_1832_),
    .A2(_2973_),
    .B(_2974_),
    .ZN(_2975_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7003_ (.A1(_2971_),
    .A2(_2975_),
    .Z(_2976_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7004_ (.A1(_1745_),
    .A2(_2967_),
    .ZN(_2977_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7005_ (.A1(_2428_),
    .A2(_2977_),
    .ZN(_2978_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7006_ (.A1(\as2650.pc[12] ),
    .A2(_2684_),
    .B1(_2978_),
    .B2(_2870_),
    .C(_2432_),
    .ZN(_2979_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7007_ (.A1(_0748_),
    .A2(_2657_),
    .B1(_2979_),
    .B2(_1939_),
    .C(_2726_),
    .ZN(_2980_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7008_ (.A1(_2976_),
    .A2(_2980_),
    .ZN(_2981_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7009_ (.A1(net38),
    .A2(_2654_),
    .B(_1461_),
    .ZN(_2982_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7010_ (.A1(_2981_),
    .A2(_2982_),
    .ZN(_0230_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7011_ (.I(net19),
    .ZN(_2983_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7012_ (.A1(_1566_),
    .A2(_1918_),
    .A3(_1635_),
    .ZN(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7013_ (.A1(_3244_),
    .A2(_1448_),
    .ZN(_2985_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7014_ (.A1(_1143_),
    .A2(_2985_),
    .B(_1620_),
    .C(_1164_),
    .ZN(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7015_ (.A1(_3140_),
    .A2(_2483_),
    .A3(_2986_),
    .ZN(_2987_));
 gf180mcu_fd_sc_mcu7t5v0__or4_1 _7016_ (.A1(_1561_),
    .A2(_2468_),
    .A3(_2984_),
    .A4(_2987_),
    .Z(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7017_ (.I(_2988_),
    .Z(_2989_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7018_ (.I(_3232_),
    .Z(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7019_ (.I(_2990_),
    .Z(_2991_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7020_ (.I(_2988_),
    .Z(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7021_ (.I(_2990_),
    .Z(_2993_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7022_ (.A1(_2993_),
    .A2(_3548_),
    .ZN(_2994_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7023_ (.A1(_3311_),
    .A2(_2991_),
    .B(_2992_),
    .C(_2994_),
    .ZN(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7024_ (.A1(_2983_),
    .A2(_2989_),
    .B(_2995_),
    .ZN(_0231_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7025_ (.I(_2990_),
    .Z(_2996_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7026_ (.I(_2990_),
    .Z(_2997_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7027_ (.A1(_2997_),
    .A2(_3529_),
    .ZN(_2998_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7028_ (.A1(_3483_),
    .A2(_2996_),
    .B(_2998_),
    .ZN(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7029_ (.I(_2988_),
    .Z(_3000_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7030_ (.A1(net30),
    .A2(_3000_),
    .ZN(_3001_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7031_ (.A1(_2989_),
    .A2(_2999_),
    .B(_3001_),
    .ZN(_0232_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7032_ (.I(_2992_),
    .Z(_3002_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7033_ (.A1(_2997_),
    .A2(_3461_),
    .ZN(_3003_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7034_ (.A1(_1710_),
    .A2(_2996_),
    .B(_3003_),
    .ZN(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7035_ (.A1(net39),
    .A2(_3000_),
    .ZN(_3005_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7036_ (.A1(_3002_),
    .A2(_3004_),
    .B(_3005_),
    .ZN(_0233_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7037_ (.A1(_2997_),
    .A2(_0976_),
    .ZN(_3006_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7038_ (.A1(_0354_),
    .A2(_2996_),
    .B(_3006_),
    .ZN(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7039_ (.A1(net40),
    .A2(_3000_),
    .ZN(_3008_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7040_ (.A1(_3002_),
    .A2(_3007_),
    .B(_3008_),
    .ZN(_0234_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7041_ (.I(net41),
    .ZN(_3009_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7042_ (.A1(_2993_),
    .A2(_0500_),
    .ZN(_3010_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7043_ (.A1(_0975_),
    .A2(_2991_),
    .B(_2992_),
    .C(_3010_),
    .ZN(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7044_ (.A1(_3009_),
    .A2(_2989_),
    .B(_3011_),
    .ZN(_0235_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7045_ (.I(net42),
    .ZN(_3012_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7046_ (.A1(_2993_),
    .A2(_0419_),
    .ZN(_3013_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7047_ (.A1(_0476_),
    .A2(_2991_),
    .B(_2988_),
    .C(_3013_),
    .ZN(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7048_ (.A1(_3012_),
    .A2(_2989_),
    .B(_3014_),
    .ZN(_0236_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7049_ (.A1(_2993_),
    .A2(_0604_),
    .ZN(_3015_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7050_ (.A1(_1728_),
    .A2(_2996_),
    .B(_3015_),
    .ZN(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7051_ (.A1(net43),
    .A2(_3000_),
    .ZN(_3017_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7052_ (.A1(_3002_),
    .A2(_3016_),
    .B(_3017_),
    .ZN(_0237_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7053_ (.A1(_0618_),
    .A2(_2997_),
    .ZN(_3018_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7054_ (.A1(_2991_),
    .A2(_2577_),
    .B(_3018_),
    .ZN(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7055_ (.A1(net44),
    .A2(_2992_),
    .ZN(_3020_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7056_ (.A1(_3002_),
    .A2(_3019_),
    .B(_3020_),
    .ZN(_0238_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7057_ (.A1(_3288_),
    .A2(_1042_),
    .ZN(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7058_ (.I(_3021_),
    .Z(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7059_ (.A1(_3287_),
    .A2(_1042_),
    .B(_3438_),
    .ZN(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7060_ (.I(_3023_),
    .Z(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7061_ (.A1(\as2650.r123[0][0] ),
    .A2(_3024_),
    .ZN(_3025_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7062_ (.A1(_3437_),
    .A2(_3022_),
    .B(_3025_),
    .ZN(_0239_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7063_ (.A1(\as2650.r123[0][1] ),
    .A2(_3024_),
    .ZN(_3026_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7064_ (.A1(_3526_),
    .A2(_3022_),
    .B(_3026_),
    .ZN(_0240_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7065_ (.A1(\as2650.r123[0][2] ),
    .A2(_3024_),
    .ZN(_3027_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7066_ (.A1(_0276_),
    .A2(_3022_),
    .B(_3027_),
    .ZN(_0241_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7067_ (.A1(\as2650.r123[0][3] ),
    .A2(_3024_),
    .ZN(_3028_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7068_ (.A1(_0365_),
    .A2(_3022_),
    .B(_3028_),
    .ZN(_0242_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7069_ (.I(_3021_),
    .Z(_3029_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7070_ (.I(_3023_),
    .Z(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7071_ (.A1(\as2650.r123[0][4] ),
    .A2(_3030_),
    .ZN(_3031_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7072_ (.A1(_0434_),
    .A2(_3029_),
    .B(_3031_),
    .ZN(_0243_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7073_ (.A1(\as2650.r123[0][5] ),
    .A2(_3030_),
    .ZN(_3032_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7074_ (.A1(_0510_),
    .A2(_3029_),
    .B(_3032_),
    .ZN(_0244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7075_ (.A1(\as2650.r123[0][6] ),
    .A2(_3030_),
    .ZN(_3033_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7076_ (.A1(_0572_),
    .A2(_3029_),
    .B(_3033_),
    .ZN(_0245_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7077_ (.A1(\as2650.r123[0][7] ),
    .A2(_3030_),
    .ZN(_3034_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7078_ (.A1(_0626_),
    .A2(_3029_),
    .B(_3034_),
    .ZN(_0246_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7079_ (.A1(_0653_),
    .A2(_1319_),
    .ZN(_3035_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7080_ (.A1(_1466_),
    .A2(_3035_),
    .ZN(_3036_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7081_ (.A1(_1544_),
    .A2(_3035_),
    .B(_3036_),
    .ZN(_0247_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7082_ (.A1(_1741_),
    .A2(_3035_),
    .ZN(_3037_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7083_ (.A1(_1234_),
    .A2(_3035_),
    .B(_3037_),
    .ZN(_0248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7084_ (.A1(_2561_),
    .A2(_1725_),
    .ZN(_3038_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7085_ (.A1(_1046_),
    .A2(_1098_),
    .B(_3038_),
    .ZN(_3039_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7086_ (.A1(_2465_),
    .A2(_0604_),
    .B(_2564_),
    .C(_1785_),
    .ZN(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7087_ (.A1(_0863_),
    .A2(_1744_),
    .A3(_0303_),
    .ZN(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7088_ (.A1(_1444_),
    .A2(_1164_),
    .A3(_1175_),
    .A4(_3041_),
    .ZN(_3042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7089_ (.A1(_1152_),
    .A2(_1178_),
    .ZN(_3043_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7090_ (.A1(_1579_),
    .A2(_1250_),
    .ZN(_3044_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7091_ (.A1(_1566_),
    .A2(_1066_),
    .B1(_1179_),
    .B2(_1173_),
    .C(_3044_),
    .ZN(_3045_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7092_ (.A1(_1137_),
    .A2(_3042_),
    .A3(_3043_),
    .A4(_3045_),
    .Z(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7093_ (.A1(_0913_),
    .A2(_0902_),
    .B(_3319_),
    .ZN(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7094_ (.A1(_2469_),
    .A2(_1165_),
    .ZN(_3048_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_1 _7095_ (.A1(_1514_),
    .A2(_2656_),
    .A3(_3047_),
    .A4(_3048_),
    .ZN(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7096_ (.A1(_3046_),
    .A2(_3049_),
    .ZN(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7097_ (.A1(_1103_),
    .A2(_1692_),
    .A3(_1150_),
    .ZN(_3051_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7098_ (.A1(_3050_),
    .A2(_3051_),
    .ZN(_3052_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7099_ (.A1(_1741_),
    .A2(_0394_),
    .B1(_3039_),
    .B2(_3040_),
    .C(_3052_),
    .ZN(_3053_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7100_ (.A1(_3050_),
    .A2(_3051_),
    .B(\as2650.psl[5] ),
    .ZN(_3054_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7101_ (.A1(_3053_),
    .A2(_3054_),
    .B(_1772_),
    .ZN(_0249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7102_ (.A1(_1046_),
    .A2(_1693_),
    .ZN(_3055_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7103_ (.A1(_1694_),
    .A2(_3055_),
    .B(_1312_),
    .ZN(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7104_ (.A1(_2465_),
    .A2(_3451_),
    .B1(_2577_),
    .B2(_1220_),
    .C(_1785_),
    .ZN(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _7105_ (.A1(_0308_),
    .A2(_0961_),
    .Z(_3058_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7106_ (.A1(_3500_),
    .A2(_3522_),
    .B(_3421_),
    .C(_3430_),
    .ZN(_3059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7107_ (.A1(_0261_),
    .A2(_0901_),
    .ZN(_3060_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7108_ (.A1(_0901_),
    .A2(_3460_),
    .B(_3060_),
    .ZN(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7109_ (.A1(_3500_),
    .A2(_3523_),
    .B1(_0273_),
    .B2(_3061_),
    .ZN(_3062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7110_ (.A1(_0274_),
    .A2(_3061_),
    .ZN(_3063_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7111_ (.A1(_3059_),
    .A2(_3062_),
    .B(_3063_),
    .ZN(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7112_ (.A1(_0308_),
    .A2(_0961_),
    .Z(_3065_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7113_ (.A1(_0445_),
    .A2(_0974_),
    .B1(_3058_),
    .B2(_3064_),
    .C(_3065_),
    .ZN(_3066_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _7114_ (.A1(_0445_),
    .A2(_0974_),
    .B1(_0466_),
    .B2(_0520_),
    .ZN(_3067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7115_ (.A1(_0466_),
    .A2(_0520_),
    .ZN(_3068_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7116_ (.A1(_0536_),
    .A2(_0581_),
    .B1(_3066_),
    .B2(_3067_),
    .C(_3068_),
    .ZN(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7117_ (.A1(_1160_),
    .A2(_0550_),
    .ZN(_3070_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7118_ (.A1(\as2650.holding_reg[7] ),
    .A2(_1160_),
    .B(_3070_),
    .ZN(_3071_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7119_ (.A1(_0537_),
    .A2(_0581_),
    .B1(_1184_),
    .B2(_3071_),
    .ZN(_3072_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7120_ (.A1(_1184_),
    .A2(_3071_),
    .ZN(_3073_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7121_ (.A1(_3069_),
    .A2(_3072_),
    .B(_3073_),
    .C(_1572_),
    .ZN(_3074_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7122_ (.A1(_1237_),
    .A2(_1692_),
    .A3(_1150_),
    .ZN(_3075_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7123_ (.A1(_3050_),
    .A2(_3075_),
    .ZN(_3076_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_1 _7124_ (.A1(_3056_),
    .A2(_3057_),
    .B(_3074_),
    .C(_3076_),
    .ZN(_3077_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7125_ (.A1(_3050_),
    .A2(_3075_),
    .B(_3411_),
    .ZN(_3078_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7126_ (.A1(_1736_),
    .A2(_3077_),
    .A3(_3078_),
    .Z(_3079_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7127_ (.I(_3079_),
    .Z(_0250_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7128_ (.A1(_3168_),
    .A2(_1711_),
    .B(_1695_),
    .ZN(_3080_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _7129_ (.A1(_0902_),
    .A2(_1177_),
    .A3(_3046_),
    .A4(_3080_),
    .Z(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__xor2_1 _7130_ (.A1(_1184_),
    .A2(_3071_),
    .Z(_3082_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7131_ (.A1(_1572_),
    .A2(_0579_),
    .ZN(_3083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7132_ (.I(_1308_),
    .Z(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7133_ (.A1(_1705_),
    .A2(_3084_),
    .B(_1834_),
    .ZN(_3085_));
 gf180mcu_fd_sc_mcu7t5v0__oai221_1 _7134_ (.A1(_3082_),
    .A2(_3083_),
    .B1(_3085_),
    .B2(_1713_),
    .C(_3081_),
    .ZN(_3086_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7135_ (.A1(\as2650.overflow ),
    .A2(_3081_),
    .B(_3086_),
    .ZN(_3087_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7136_ (.A1(_1772_),
    .A2(_3087_),
    .ZN(_0251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7137_ (.A1(_1720_),
    .A2(_1567_),
    .ZN(_3088_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7138_ (.A1(_1301_),
    .A2(_1065_),
    .ZN(_3089_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7139_ (.A1(_1071_),
    .A2(_1087_),
    .A3(_3089_),
    .ZN(_3090_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7140_ (.A1(_1056_),
    .A2(_1108_),
    .B(_3090_),
    .ZN(_3091_));
 gf180mcu_fd_sc_mcu7t5v0__oai31_1 _7141_ (.A1(_1076_),
    .A2(_1118_),
    .A3(_1086_),
    .B(_3091_),
    .ZN(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7142_ (.A1(_3088_),
    .A2(_3092_),
    .ZN(_3093_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7143_ (.A1(_3432_),
    .A2(_3093_),
    .ZN(_3094_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7144_ (.A1(_1720_),
    .A2(_1703_),
    .A3(_3084_),
    .ZN(_3095_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7145_ (.A1(_1722_),
    .A2(_3093_),
    .A3(_3095_),
    .Z(_3096_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7146_ (.A1(_2496_),
    .A2(_3094_),
    .A3(_3096_),
    .ZN(_0252_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7147_ (.A1(_1715_),
    .A2(_1567_),
    .ZN(_3097_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7148_ (.A1(_3092_),
    .A2(_3097_),
    .ZN(_3098_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7149_ (.A1(_3319_),
    .A2(_3098_),
    .ZN(_3099_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7150_ (.A1(_1715_),
    .A2(_1703_),
    .A3(_3084_),
    .ZN(_3100_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7151_ (.A1(_1717_),
    .A2(_3098_),
    .A3(_3100_),
    .Z(_3101_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7152_ (.A1(_2496_),
    .A2(_3099_),
    .A3(_3101_),
    .ZN(_0253_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7153_ (.A1(_1333_),
    .A2(_1692_),
    .ZN(_3102_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7154_ (.A1(_3092_),
    .A2(_3102_),
    .ZN(_3103_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7155_ (.A1(\as2650.psl[1] ),
    .A2(_3103_),
    .ZN(_3104_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7156_ (.A1(_1333_),
    .A2(_1703_),
    .A3(_3084_),
    .ZN(_3105_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _7157_ (.A1(_1706_),
    .A2(_3103_),
    .A3(_3105_),
    .Z(_3106_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7158_ (.A1(_1116_),
    .A2(_3104_),
    .A3(_3106_),
    .ZN(_0254_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _7159_ (.A1(_1651_),
    .A2(_1131_),
    .B(_1072_),
    .C(_1087_),
    .ZN(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _7160_ (.I(_3107_),
    .ZN(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7161_ (.A1(_1349_),
    .A2(_1733_),
    .B(_3108_),
    .ZN(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7162_ (.A1(_1105_),
    .A2(_1109_),
    .ZN(_3110_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _7163_ (.A1(_1728_),
    .A2(_1729_),
    .B1(_3110_),
    .B2(_1236_),
    .ZN(_3111_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _7164_ (.A1(_1290_),
    .A2(_3109_),
    .B1(_3111_),
    .B2(_3108_),
    .C(_1595_),
    .ZN(_0255_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7165_ (.I(_3107_),
    .Z(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7166_ (.A1(_3088_),
    .A2(_3112_),
    .Z(_3113_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7167_ (.I(_1109_),
    .Z(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7168_ (.A1(_3114_),
    .A2(_1721_),
    .B(_1722_),
    .ZN(_3115_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7169_ (.A1(_3113_),
    .A2(_3115_),
    .ZN(_3116_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7170_ (.A1(_1288_),
    .A2(_3113_),
    .B(_3116_),
    .C(_1691_),
    .ZN(_0256_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _7171_ (.A1(_3097_),
    .A2(_3107_),
    .Z(_3117_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7172_ (.A1(_3114_),
    .A2(_1716_),
    .B(_1717_),
    .ZN(_3118_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7173_ (.A1(_3117_),
    .A2(_3118_),
    .ZN(_3119_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _7174_ (.A1(_2533_),
    .A2(_3117_),
    .B(_3119_),
    .C(_1798_),
    .ZN(_0257_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7175_ (.A1(_1711_),
    .A2(_3112_),
    .ZN(_3120_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7176_ (.A1(_1710_),
    .A2(_1729_),
    .B(_3110_),
    .ZN(_3121_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7177_ (.A1(\as2650.psu[2] ),
    .A2(_3120_),
    .B(_1460_),
    .ZN(_3122_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7178_ (.A1(_3120_),
    .A2(_3121_),
    .B(_3122_),
    .ZN(_0258_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7179_ (.A1(_3114_),
    .A2(_1704_),
    .B(_1706_),
    .ZN(_3123_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _7180_ (.A1(_3102_),
    .A2(_3112_),
    .A3(_3123_),
    .ZN(_3124_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7181_ (.A1(_3102_),
    .A2(_3112_),
    .ZN(_3125_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7182_ (.A1(\as2650.psu[1] ),
    .A2(_3125_),
    .B(_1461_),
    .ZN(_3126_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _7183_ (.A1(_3124_),
    .A2(_3126_),
    .ZN(_0259_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_1 _7184_ (.A1(_1237_),
    .A2(_1733_),
    .B(_3108_),
    .ZN(_3127_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7185_ (.A1(\as2650.psu[0] ),
    .A2(_3127_),
    .ZN(_3128_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _7186_ (.A1(_3114_),
    .A2(_1693_),
    .ZN(_3129_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _7187_ (.A1(_1694_),
    .A2(_3108_),
    .A3(_3129_),
    .ZN(_3130_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _7188_ (.A1(_3128_),
    .A2(_3130_),
    .B(_2496_),
    .ZN(_0260_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7189_ (.D(_0000_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7190_ (.D(_0001_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7191_ (.D(_0002_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7192_ (.D(_0003_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7193_ (.D(_0004_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7194_ (.D(_0005_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7195_ (.D(_0006_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7196_ (.D(_0007_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.r123[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7197_ (.D(_0008_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7198_ (.D(_0009_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7199_ (.D(_0010_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7200_ (.D(_0011_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7201_ (.D(_0012_),
    .CLK(clknet_leaf_61_wb_clk_i),
    .Q(\as2650.r123[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7202_ (.D(_0013_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7203_ (.D(_0014_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7204_ (.D(_0015_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7205_ (.D(_0016_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7206_ (.D(_0017_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7207_ (.D(_0018_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7208_ (.D(_0019_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[4][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7209_ (.D(_0020_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7210_ (.D(_0021_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7211_ (.D(_0022_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7212_ (.D(_0023_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7213_ (.D(_0024_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[4][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7214_ (.D(_0025_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7215_ (.D(_0026_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7216_ (.D(_0027_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[4][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7217_ (.D(_0028_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[4][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7218_ (.D(_0029_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7219_ (.D(_0030_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7220_ (.D(_0031_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7221_ (.D(_0032_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7222_ (.D(_0033_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7223_ (.D(_0034_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7224_ (.D(_0035_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7225_ (.D(_0036_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7226_ (.D(_0037_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[3][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7227_ (.D(_0038_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7228_ (.D(_0039_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7229_ (.D(_0040_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7230_ (.D(_0041_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7231_ (.D(_0042_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7232_ (.D(_0043_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7233_ (.D(_0044_),
    .CLK(clknet_leaf_24_wb_clk_i),
    .Q(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7234_ (.D(_0045_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7235_ (.D(_0046_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7236_ (.D(_0047_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7237_ (.D(_0048_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7238_ (.D(_0049_),
    .CLK(clknet_leaf_36_wb_clk_i),
    .Q(\as2650.stack[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7239_ (.D(_0050_),
    .CLK(clknet_leaf_39_wb_clk_i),
    .Q(\as2650.stack[2][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7240_ (.D(_0051_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7241_ (.D(_0052_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7242_ (.D(_0053_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7243_ (.D(_0054_),
    .CLK(clknet_leaf_31_wb_clk_i),
    .Q(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7244_ (.D(_0055_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7245_ (.D(_0056_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7246_ (.D(_0057_),
    .CLK(clknet_leaf_48_wb_clk_i),
    .Q(\as2650.stack[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7247_ (.D(_0058_),
    .CLK(clknet_leaf_46_wb_clk_i),
    .Q(\as2650.stack[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7248_ (.D(_0059_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7249_ (.D(_0060_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7250_ (.D(_0061_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7251_ (.D(_0062_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7252_ (.D(_0063_),
    .CLK(clknet_leaf_41_wb_clk_i),
    .Q(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7253_ (.D(_0064_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[1][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7254_ (.D(_0065_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[1][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7255_ (.D(_0066_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7256_ (.D(_0067_),
    .CLK(clknet_leaf_38_wb_clk_i),
    .Q(\as2650.stack[1][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7257_ (.D(_0068_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7258_ (.D(_0069_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7259_ (.D(_0070_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7260_ (.D(_0071_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7261_ (.D(_0072_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7262_ (.D(_0073_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7263_ (.D(_0074_),
    .CLK(clknet_leaf_40_wb_clk_i),
    .Q(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7264_ (.D(_0075_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7265_ (.D(_0076_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7266_ (.D(_0077_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[0][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7267_ (.D(_0078_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[0][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7268_ (.D(_0079_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[0][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7269_ (.D(_0080_),
    .CLK(clknet_leaf_32_wb_clk_i),
    .Q(\as2650.stack[0][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7270_ (.D(_0081_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7271_ (.D(_0082_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7272_ (.D(_0083_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7273_ (.D(_0084_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7274_ (.D(_0085_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123_2[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7275_ (.D(_0086_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7276_ (.D(_0087_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[2][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7277_ (.D(_0088_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r123_2[2][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7278_ (.D(_0089_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.psu[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7279_ (.D(_0090_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.psl[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7280_ (.D(_0091_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.psl[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7281_ (.D(_0092_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7282_ (.D(_0093_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7283_ (.D(_0094_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.ins_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7284_ (.D(_0095_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7285_ (.D(_0096_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7286_ (.D(_0097_),
    .CLK(clknet_leaf_8_wb_clk_i),
    .Q(\as2650.ins_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7287_ (.D(_0098_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7288_ (.D(_0099_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7289_ (.D(_0100_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[6][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7290_ (.D(_0101_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[6][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7291_ (.D(_0102_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7292_ (.D(_0103_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7293_ (.D(_0104_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7294_ (.D(_0105_),
    .CLK(clknet_leaf_43_wb_clk_i),
    .Q(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7295_ (.D(_0106_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[6][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7296_ (.D(_0107_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7297_ (.D(_0108_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7298_ (.D(_0109_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7299_ (.D(_0110_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[6][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7300_ (.D(_0111_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123_2[1][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7301_ (.D(_0112_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[1][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7302_ (.D(_0113_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7303_ (.D(_0114_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7304_ (.D(_0115_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7305_ (.D(_0116_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7306_ (.D(_0117_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7307_ (.D(_0118_),
    .CLK(clknet_leaf_62_wb_clk_i),
    .Q(\as2650.r123_2[1][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7308_ (.D(_0119_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.r123[3][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7309_ (.D(_0120_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7310_ (.D(_0121_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7311_ (.D(_0122_),
    .CLK(clknet_leaf_56_wb_clk_i),
    .Q(\as2650.r123[3][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7312_ (.D(_0123_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7313_ (.D(_0124_),
    .CLK(clknet_leaf_55_wb_clk_i),
    .Q(\as2650.r123[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7314_ (.D(_0125_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.r123[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7315_ (.D(_0126_),
    .CLK(clknet_leaf_57_wb_clk_i),
    .Q(\as2650.r123[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7316_ (.D(_0127_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7317_ (.D(_0128_),
    .CLK(clknet_leaf_50_wb_clk_i),
    .Q(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7318_ (.D(_0129_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[5][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7319_ (.D(_0130_),
    .CLK(clknet_leaf_51_wb_clk_i),
    .Q(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7320_ (.D(_0131_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7321_ (.D(_0132_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7322_ (.D(_0133_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7323_ (.D(_0134_),
    .CLK(clknet_leaf_42_wb_clk_i),
    .Q(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7324_ (.D(_0135_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[5][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7325_ (.D(_0136_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7326_ (.D(_0137_),
    .CLK(clknet_leaf_37_wb_clk_i),
    .Q(\as2650.stack[5][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7327_ (.D(_0138_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7328_ (.D(_0139_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[5][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7329_ (.D(_0140_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7330_ (.D(_0141_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7331_ (.D(_0142_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7332_ (.D(_0143_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123_2[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7333_ (.D(_0144_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7334_ (.D(_0145_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7335_ (.D(_0146_),
    .CLK(clknet_leaf_64_wb_clk_i),
    .Q(\as2650.r123_2[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7336_ (.D(_0147_),
    .CLK(clknet_leaf_1_wb_clk_i),
    .Q(\as2650.r123_2[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7337_ (.D(_0148_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7338_ (.D(_0149_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7339_ (.D(_0150_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123_2[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7340_ (.D(_0151_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7341_ (.D(_0152_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7342_ (.D(_0153_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7343_ (.D(_0154_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7344_ (.D(_0155_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7345_ (.D(_0156_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7346_ (.D(_0157_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7347_ (.D(_0158_),
    .CLK(clknet_leaf_13_wb_clk_i),
    .Q(\as2650.addr_buff[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7348_ (.D(_0159_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(net21));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7349_ (.D(_0160_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7350_ (.D(_0161_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(net20));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7351_ (.D(_0162_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(net23));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7352_ (.D(_0163_),
    .CLK(clknet_leaf_21_wb_clk_i),
    .Q(net22));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7353_ (.D(_0164_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.idx_ctrl[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7354_ (.D(_0165_),
    .CLK(clknet_leaf_12_wb_clk_i),
    .Q(\as2650.idx_ctrl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7355_ (.D(_0166_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7356_ (.D(_0167_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.holding_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7357_ (.D(_0168_),
    .CLK(clknet_leaf_65_wb_clk_i),
    .Q(\as2650.holding_reg[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7358_ (.D(_0169_),
    .CLK(clknet_3_0_0_wb_clk_i),
    .Q(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7359_ (.D(_0170_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7360_ (.D(_0171_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.holding_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7361_ (.D(_0172_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7362_ (.D(_0173_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7363_ (.D(_0174_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7364_ (.D(_0175_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.cycle[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7365_ (.D(_0176_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.cycle[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7366_ (.D(_0177_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(\as2650.cycle[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7367_ (.D(_0178_),
    .CLK(clknet_leaf_16_wb_clk_i),
    .Q(\as2650.cycle[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7368_ (.D(_0179_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7369_ (.D(_0180_),
    .CLK(clknet_leaf_17_wb_clk_i),
    .Q(\as2650.cycle[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7370_ (.D(_0181_),
    .CLK(clknet_leaf_19_wb_clk_i),
    .Q(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7371_ (.D(_0182_),
    .CLK(clknet_3_3_0_wb_clk_i),
    .Q(\as2650.cycle[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7372_ (.D(_0183_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.psu[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7373_ (.D(_0184_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7374_ (.D(_0185_),
    .CLK(clknet_3_5_0_wb_clk_i),
    .Q(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7375_ (.D(_0186_),
    .CLK(clknet_leaf_47_wb_clk_i),
    .Q(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7376_ (.D(_0187_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7377_ (.D(_0188_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7378_ (.D(_0189_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7379_ (.D(_0190_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7380_ (.D(_0191_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7381_ (.D(_0192_),
    .CLK(clknet_leaf_30_wb_clk_i),
    .Q(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7382_ (.D(_0193_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7383_ (.D(_0194_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7384_ (.D(_0195_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.pc[11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7385_ (.D(_0196_),
    .CLK(clknet_leaf_25_wb_clk_i),
    .Q(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7386_ (.D(_0197_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7387_ (.D(_0198_),
    .CLK(clknet_3_1_0_wb_clk_i),
    .Q(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7388_ (.D(_0199_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7389_ (.D(_0200_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7390_ (.D(_0201_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7391_ (.D(_0202_),
    .CLK(clknet_leaf_10_wb_clk_i),
    .Q(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7392_ (.D(_0203_),
    .CLK(clknet_leaf_9_wb_clk_i),
    .Q(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7393_ (.D(_0204_),
    .CLK(clknet_3_2_0_wb_clk_i),
    .Q(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7394_ (.D(_0205_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7395_ (.D(_0206_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7396_ (.D(_0207_),
    .CLK(clknet_leaf_49_wb_clk_i),
    .Q(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7397_ (.D(_0208_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7398_ (.D(_0209_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7399_ (.D(_0210_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7400_ (.D(_0211_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7401_ (.D(_0212_),
    .CLK(clknet_leaf_45_wb_clk_i),
    .Q(\as2650.stack[7][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7402_ (.D(_0213_),
    .CLK(clknet_leaf_44_wb_clk_i),
    .Q(\as2650.stack[7][8] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7403_ (.D(_0214_),
    .CLK(clknet_leaf_35_wb_clk_i),
    .Q(\as2650.stack[7][9] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7404_ (.D(_0215_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][10] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7405_ (.D(_0216_),
    .CLK(clknet_leaf_34_wb_clk_i),
    .Q(\as2650.stack[7][11] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7406_ (.D(_0217_),
    .CLK(clknet_leaf_33_wb_clk_i),
    .Q(\as2650.stack[7][12] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7407_ (.D(_0218_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net25));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7408_ (.D(_0219_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net26));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7409_ (.D(_0220_),
    .CLK(clknet_opt_3_1_wb_clk_i),
    .Q(net27));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7410_ (.D(_0221_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net28));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7411_ (.D(_0222_),
    .CLK(clknet_leaf_27_wb_clk_i),
    .Q(net29));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7412_ (.D(_0223_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net31));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7413_ (.D(_0224_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net32));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7414_ (.D(_0225_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net33));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7415_ (.D(_0226_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net34));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7416_ (.D(_0227_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net35));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7417_ (.D(_0228_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net36));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7418_ (.D(_0229_),
    .CLK(clknet_leaf_29_wb_clk_i),
    .Q(net37));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7419_ (.D(_0230_),
    .CLK(clknet_leaf_28_wb_clk_i),
    .Q(net38));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7420_ (.D(_0231_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net19));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7421_ (.D(_0232_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net30));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7422_ (.D(_0233_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net39));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7423_ (.D(_0234_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net40));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7424_ (.D(_0235_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net41));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7425_ (.D(_0236_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net42));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7426_ (.D(_0237_),
    .CLK(clknet_leaf_15_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7427_ (.D(_0238_),
    .CLK(clknet_leaf_14_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7428_ (.D(_0239_),
    .CLK(clknet_leaf_2_wb_clk_i),
    .Q(\as2650.r123[0][0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7429_ (.D(_0240_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[0][1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7430_ (.D(_0241_),
    .CLK(clknet_leaf_0_wb_clk_i),
    .Q(\as2650.r123[0][2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7431_ (.D(_0242_),
    .CLK(clknet_leaf_63_wb_clk_i),
    .Q(\as2650.r123[0][3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7432_ (.D(_0243_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[0][4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7433_ (.D(_0244_),
    .CLK(clknet_leaf_3_wb_clk_i),
    .Q(\as2650.r123[0][5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7434_ (.D(_0245_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7435_ (.D(_0246_),
    .CLK(clknet_leaf_4_wb_clk_i),
    .Q(\as2650.r123[0][7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7436_ (.D(_0247_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.ins_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7437_ (.D(_0248_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7438_ (.D(_0249_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7439_ (.D(_0250_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7440_ (.D(_0251_),
    .CLK(clknet_leaf_6_wb_clk_i),
    .Q(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _7441_ (.D(_0252_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7442_ (.D(_0253_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7443_ (.D(_0254_),
    .CLK(clknet_3_4_0_wb_clk_i),
    .Q(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7444_ (.D(_0255_),
    .CLK(clknet_leaf_52_wb_clk_i),
    .Q(net24));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7445_ (.D(_0256_),
    .CLK(clknet_leaf_60_wb_clk_i),
    .Q(\as2650.psu[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7446_ (.D(_0257_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7447_ (.D(_0258_),
    .CLK(clknet_leaf_53_wb_clk_i),
    .Q(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7448_ (.D(_0259_),
    .CLK(clknet_leaf_54_wb_clk_i),
    .Q(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _7449_ (.D(_0260_),
    .CLK(clknet_leaf_7_wb_clk_i),
    .Q(\as2650.psu[0] ));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_0_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_54 (.ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_55 (.ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_56 (.ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_57 (.ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_58 (.ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_59 (.ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_60 (.ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_61 (.ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_62 (.ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_63 (.ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_64 (.ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_65 (.ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_66 (.ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_67 (.ZN(net67));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_68 (.ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_69 (.ZN(net69));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_70 (.ZN(net70));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_71 (.ZN(net71));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_72 (.ZN(net72));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_73 (.ZN(net73));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_74 (.ZN(net74));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_75 (.ZN(net75));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_76 (.ZN(net76));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_77 (.ZN(net77));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_78 (.ZN(net78));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_79 (.ZN(net79));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_80 (.ZN(net80));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_81 (.ZN(net81));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_82 (.ZN(net82));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_83 (.ZN(net83));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_84 (.ZN(net84));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_85 (.ZN(net85));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_86 (.ZN(net86));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_87 (.ZN(net87));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_88 (.ZN(net88));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_89 (.ZN(net89));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_90 (.ZN(net90));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_91 (.ZN(net91));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_92 (.ZN(net92));
 gf180mcu_fd_sc_mcu7t5v0__tieh wrapped_as2650_93 (.Z(net93));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7491_ (.I(net46),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7492_ (.I(net46),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7493_ (.I(net47),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7494_ (.I(net47),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7495_ (.I(net47),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7496_ (.I(net46),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _7497_ (.I(net46),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_9 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_110 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_111 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_112 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_113 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_114 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_115 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_116 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_117 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_118 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_119 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_120 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_121 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_122 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_123 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_124 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_125 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_126 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_127 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_128 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_129 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_130 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_131 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_132 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_133 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_134 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_135 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_136 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_137 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_138 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_139 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_140 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_141 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_142 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_143 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_144 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_145 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_146 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_147 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_148 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_149 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_150 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_151 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_152 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_153 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_154 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_155 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_156 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_157 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_158 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_159 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_160 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_161 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_162 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_163 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_164 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_165 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_166 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_167 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_168 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_169 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_170 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_171 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_172 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_173 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_174 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_175 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_176 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_177 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_178 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_179 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_180 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_181 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_182 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_183 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_184 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_185 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_186 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_187 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_188 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_189 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_190 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_191 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_192 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_193 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_194 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_195 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_196 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_197 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_198 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_199 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_200 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_201 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_202 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_203 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_204 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_205 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_206 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_207 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_208 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_209 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_210 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_211 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_212 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_213 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_214 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_215 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_216 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_217 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_218 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_219 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_220 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_221 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_222 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_223 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_224 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_225 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_226 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_227 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_228 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_229 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_230 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_231 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_232 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_233 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_234 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_235 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_236 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_237 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_238 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_239 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_240 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_241 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_242 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_243 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_244 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_245 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_246 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_247 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_248 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_249 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_250 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_251 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_252 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_253 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_254 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_255 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_256 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_257 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_258 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_259 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_260 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_261 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_262 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_263 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_264 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_265 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_266 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_267 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_268 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_269 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_270 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_271 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_272 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_273 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_274 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_275 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_276 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_277 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_278 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_279 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_280 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_281 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_282 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_283 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_284 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_285 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_286 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_287 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_288 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_1999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2525 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2526 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2527 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2528 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2529 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2530 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2531 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2532 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2533 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2534 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2535 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2536 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2537 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2538 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2539 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2540 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2541 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2542 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2543 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2544 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2545 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2546 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2547 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2548 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2549 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2550 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2551 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2552 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2553 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2554 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2555 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2556 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2557 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2558 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2559 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2560 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2561 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2562 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2563 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2564 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2565 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2566 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2567 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2568 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2569 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2570 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2571 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2572 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2573 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2574 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2575 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2576 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2577 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2578 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2579 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2580 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2581 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2582 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2583 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2584 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2585 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2586 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2587 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2588 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2589 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2590 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2591 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2592 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2593 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2594 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2595 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2596 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2597 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2598 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2599 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2600 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2601 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2602 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2603 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2604 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2605 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2606 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2607 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2608 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2609 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2610 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2611 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2612 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2613 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2614 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2615 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2616 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2617 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2618 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2619 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2620 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2621 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2622 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2623 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2624 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2625 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2626 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2627 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2628 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2629 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2630 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2631 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2632 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2633 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2634 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2635 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2636 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2637 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2638 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2639 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2640 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2641 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2642 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2643 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2644 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2645 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2646 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2647 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2648 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2649 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2650 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2651 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2652 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2653 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2654 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2655 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2656 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2657 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2658 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2659 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2660 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2661 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2662 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2663 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2664 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2665 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2666 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2667 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2668 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2669 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2670 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2671 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2672 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2673 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2674 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2675 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2676 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2677 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2678 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2679 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2680 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2681 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2682 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2683 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2684 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2685 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2686 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2687 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2688 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2689 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2690 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2691 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2692 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2693 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2694 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2695 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2696 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2697 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2698 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2699 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2700 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2701 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2702 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2703 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2704 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2705 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2706 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2707 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2708 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2709 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2710 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2711 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2712 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2713 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2714 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2715 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2716 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2717 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2718 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2719 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2720 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2721 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2722 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2723 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2724 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2725 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2726 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2727 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2728 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2729 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2730 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2731 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2732 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2733 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2734 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2735 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2736 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2737 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2738 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2739 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2740 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2741 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2742 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2743 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2744 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2745 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2746 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2747 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2748 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2749 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2750 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2751 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2752 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2753 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2754 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2755 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2756 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2757 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2758 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2759 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2760 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2761 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2762 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2763 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2764 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2765 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2766 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2767 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2768 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2769 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2770 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2771 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2772 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2773 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2774 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2775 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2776 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2777 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2778 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2779 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2780 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2781 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2782 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2783 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2784 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2785 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2786 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2787 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2788 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2789 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2790 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2791 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2792 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2793 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2794 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2795 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2796 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2797 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2798 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2799 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2800 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2801 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2802 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2803 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2804 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2805 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2806 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2807 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2808 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2809 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2810 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2811 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2812 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2813 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2814 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2815 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2816 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2817 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2818 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2819 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2820 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2821 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2822 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2823 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2824 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2825 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2826 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2827 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2828 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2829 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2830 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2831 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2832 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2833 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2834 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2835 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2836 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2837 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2838 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2839 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2840 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2841 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2842 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2843 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2844 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2845 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2846 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2847 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2848 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2849 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2850 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2851 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2852 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2853 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2854 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2855 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2856 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2857 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2858 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2859 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2860 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2861 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2862 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2863 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2864 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2865 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2866 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2867 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2868 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2869 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2870 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2871 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2872 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2873 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2874 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2875 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2876 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2877 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2878 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2879 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2880 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2881 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2882 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2883 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2884 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2885 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2886 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2887 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2888 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2889 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2890 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2891 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2892 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2893 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2894 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2895 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2896 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2897 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2898 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2899 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2900 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2901 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2902 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2903 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2904 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2905 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2906 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2907 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2908 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2909 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2910 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2911 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2912 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2913 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2914 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2915 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2916 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2917 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2918 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2919 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2920 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2921 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2922 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2923 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2924 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2925 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2926 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2927 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2928 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2929 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2930 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2931 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2932 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2933 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2934 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2935 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2936 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2937 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2938 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2939 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2940 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2941 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2942 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2943 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2944 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2945 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2946 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2947 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2948 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2949 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2950 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2951 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2952 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2953 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2954 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2955 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2956 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2957 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2958 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2959 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2960 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2961 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2962 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2963 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2964 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2965 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2966 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2967 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2968 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2969 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2970 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2971 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2972 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2973 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2974 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2975 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2976 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2977 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2978 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2979 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2980 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2981 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2982 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2983 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2984 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2985 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2986 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2987 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2988 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2989 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2990 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2991 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2992 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2993 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2994 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2995 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2996 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2997 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2998 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_2999 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3000 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3001 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3002 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3003 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3004 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3005 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3006 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3007 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3008 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3009 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3010 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3011 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3012 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3013 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3014 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3015 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3016 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3017 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3018 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3019 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3020 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3021 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3022 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3023 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3024 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3025 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3026 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3027 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3028 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3029 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3030 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3031 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3032 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3033 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3034 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3035 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3036 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3037 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3038 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3039 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3040 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3041 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3042 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3043 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3044 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3045 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3046 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3047 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3048 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3049 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3050 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3051 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3052 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3053 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3054 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3055 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3056 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3057 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3058 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3059 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3060 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3061 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3062 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3063 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3064 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3065 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3066 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3067 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3068 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3069 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3070 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3071 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3072 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3073 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3074 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3075 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3076 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3077 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3078 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3079 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3080 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3081 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3082 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3083 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3084 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3085 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3086 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3087 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3088 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3089 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3090 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3091 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3092 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3093 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3094 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3095 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3096 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3097 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3098 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3099 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3100 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3101 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3102 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3103 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3104 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3105 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3106 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3107 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3108 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3109 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3170 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3425 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3426 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3427 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3428 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3429 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3430 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3431 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3432 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3433 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3434 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3435 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3436 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3437 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3438 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3439 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3440 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3441 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3442 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3443 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3444 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3445 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3446 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3447 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3448 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3449 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3450 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3451 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3452 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3453 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3454 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3455 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3456 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3457 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3458 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3459 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3460 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3461 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3462 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3463 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3464 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3465 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3466 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3467 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3468 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3469 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3470 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3471 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3472 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3473 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3474 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3475 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3476 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3477 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3478 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3479 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3480 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3481 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3482 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3483 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3484 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3485 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3486 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3487 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3488 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3489 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3490 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3491 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3492 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3493 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3494 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3495 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3496 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3497 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3498 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3499 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3500 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3501 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3502 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3503 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3504 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3505 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3506 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3507 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3508 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3509 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3510 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3511 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3512 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3513 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3514 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3515 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3516 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3517 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3518 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3519 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3520 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3521 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3522 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3523 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3524 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_3525 ();
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(io_in[0]),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input2 (.I(io_in[1]),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input3 (.I(io_in[2]),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input4 (.I(io_in[3]),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input5 (.I(io_in[4]),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input6 (.I(io_in[5]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 input7 (.I(io_in[6]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input8 (.I(io_in[7]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 input9 (.I(io_in[8]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input10 (.I(wb_rst_i),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output11 (.I(net11),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output12 (.I(net12),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output13 (.I(net13),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output14 (.I(net14),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output15 (.I(net15),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output16 (.I(net16),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output17 (.I(net17),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output18 (.I(net49),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output19 (.I(net19),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output20 (.I(net20),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output21 (.I(net21),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output22 (.I(net22),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output23 (.I(net23),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output24 (.I(net24),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output25 (.I(net25),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output26 (.I(net52),
    .Z(io_out[16]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output27 (.I(net27),
    .Z(io_out[17]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output28 (.I(net28),
    .Z(io_out[18]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output29 (.I(net29),
    .Z(io_out[19]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output30 (.I(net30),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output31 (.I(net31),
    .Z(io_out[20]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output32 (.I(net32),
    .Z(io_out[21]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output33 (.I(net33),
    .Z(io_out[22]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output34 (.I(net34),
    .Z(io_out[23]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output35 (.I(net35),
    .Z(io_out[24]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output36 (.I(net36),
    .Z(io_out[25]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output37 (.I(net37),
    .Z(io_out[26]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output38 (.I(net38),
    .Z(io_out[27]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output39 (.I(net39),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output40 (.I(net40),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output41 (.I(net41),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output42 (.I(net42),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output43 (.I(net43),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output44 (.I(net44),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 output45 (.I(net45),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__dlyc_1 fanout46 (.I(net48),
    .Z(net46));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout47 (.I(net48),
    .Z(net47));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout48 (.I(net49),
    .Z(net48));
 gf180mcu_fd_sc_mcu7t5v0__dlyb_1 fanout49 (.I(net18),
    .Z(net49));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout50 (.I(net34),
    .Z(net50));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 fanout51 (.I(net31),
    .Z(net51));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 fanout52 (.I(net26),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__tiel wrapped_as2650_53 (.ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_1_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_2_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_3_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_4_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_4_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_6_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_7_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_8_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_8_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_9_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_9_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_10_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_10_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_12_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_12_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_13_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_13_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_14_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_15_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_16_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_16_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_17_wb_clk_i (.I(clknet_3_2_0_wb_clk_i),
    .Z(clknet_leaf_17_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_19_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_21_wb_clk_i (.I(clknet_opt_1_0_wb_clk_i),
    .Z(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_24_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_24_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_25_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_27_wb_clk_i (.I(clknet_opt_4_0_wb_clk_i),
    .Z(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_28_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_28_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_29_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_30_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_30_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_31_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_32_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_33_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_34_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_35_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_36_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_37_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_38_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_39_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_40_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_41_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_41_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_42_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_43_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_43_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_44_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_45_wb_clk_i (.I(clknet_3_7_0_wb_clk_i),
    .Z(clknet_leaf_45_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_46_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_46_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_47_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_leaf_47_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_48_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_49_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_50_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_51_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_51_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_52_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_53_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_54_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_55_wb_clk_i (.I(clknet_opt_2_1_wb_clk_i),
    .Z(clknet_leaf_55_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_56_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_56_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_57_wb_clk_i (.I(clknet_3_4_0_wb_clk_i),
    .Z(clknet_leaf_57_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_60_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_61_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_61_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_62_wb_clk_i (.I(clknet_3_1_0_wb_clk_i),
    .Z(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_63_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_63_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_64_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_leaf_65_wb_clk_i (.I(clknet_3_0_0_wb_clk_i),
    .Z(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_0_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_1_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_2_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_3_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_4_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_5_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_6_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 clkbuf_3_7_0_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_1_0_wb_clk_i (.I(clknet_3_3_0_wb_clk_i),
    .Z(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_0_wb_clk_i (.I(clknet_3_5_0_wb_clk_i),
    .Z(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_2_1_wb_clk_i (.I(clknet_opt_2_0_wb_clk_i),
    .Z(clknet_opt_2_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_3_1_wb_clk_i (.I(clknet_opt_3_0_wb_clk_i),
    .Z(clknet_opt_3_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_opt_4_0_wb_clk_i (.I(clknet_3_6_0_wb_clk_i),
    .Z(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__D (.I(_0093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__D (.I(_0094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7345__D (.I(_0156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7353__D (.I(_0164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7354__D (.I(_0165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7364__D (.I(_0175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7365__D (.I(_0176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__D (.I(_0177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7367__D (.I(_0178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__D (.I(_0182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7377__D (.I(_0188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__D (.I(_0195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__D (.I(_0197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__D (.I(_0199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7389__D (.I(_0200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7390__D (.I(_0201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7391__D (.I(_0202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7392__D (.I(_0203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__D (.I(_0204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A3 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A1 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4063__A2 (.I(_0263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4098__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A2 (.I(_0265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6510__A1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4072__B1 (.I(_0268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A2 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4191__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4070__A1 (.I(_0269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A3 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__A1 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A2 (.I(_0274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4917__I (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A2 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A1 (.I(_0278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__C (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4194__S (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A1 (.I(_0279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A1 (.I(_0281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4106__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4083__I (.I(_0282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A3 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A4 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A3 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4084__A2 (.I(_0283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4115__A2 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4096__A3 (.I(_0285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4186__B (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A2 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4087__A1 (.I(_0286_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5078__B (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A2 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4099__B (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4091__A1 (.I(_0288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__A1 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__A1 (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__C (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4101__B (.I(_0300_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A3 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__B2 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A1 (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__C (.I(_0303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B2 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A1 (.I(_0305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A4 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__B (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4117__I (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4108__A2 (.I(_0306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A1 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4177__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4109__A2 (.I(_0308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A1 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__C (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4111__B2 (.I(_0310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A2 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4264__C (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4193__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4113__A1 (.I(_0312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A2 (.I(_0315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4222__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4146__I (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4130__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__A2 (.I(_0317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__B2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__A1 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4124__B2 (.I(_0319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A1 (.I(_0320_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4129__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4123__A2 (.I(_0321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6783__A2 (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4125__I (.I(_0324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4852__A1 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4126__A2 (.I(_0325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6791__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6789__A2 (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4131__I (.I(_0330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4850__A1 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__A2 (.I(_0331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__B2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__B1 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4153__A2 (.I(_0332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4288__S (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4216__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4213__A1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__S1 (.I(_0333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A1 (.I(_0335_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5060__I (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A1 (.I(_0336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__A2 (.I(_0337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4170__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4140__A2 (.I(_0339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A4 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4199__A1 (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4141__I (.I(_0340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__C2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A2 (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4142__I (.I(_0341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4846__A1 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4302__I (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4152__A2 (.I(_0342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6782__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A1 (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4144__I (.I(_0343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6755__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__B1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A1 (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4145__I (.I(_0344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5129__I (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4844__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4151__A1 (.I(_0345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__A2 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4858__I (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4149__A1 (.I(_0346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4845__A1 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4150__A2 (.I(_0349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7038__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A1 (.I(_0354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5041__I (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5011__I (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4918__I (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4156__I (.I(_0355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A1 (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4157__I (.I(_0356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A2 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4990__I (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A1 (.I(_0357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A2 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4778__A1 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A3 (.I(_0358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4160__A2 (.I(_0359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A1 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A2 (.I(_0365_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4173__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4171__I (.I(_0369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4204__I (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4172__A2 (.I(_0370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A3 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4279__I (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4174__A2 (.I(_0372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4179__A2 (.I(_0377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5047__I (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4182__A1 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4181__A2 (.I(_0379_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__C (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4333__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4245__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__A1 (.I(_0383_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A1 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A2 (.I(_0394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4270__A1 (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4197__I (.I(_0395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A2 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4198__A1 (.I(_0396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A2 (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4201__I (.I(_0399_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6542__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4868__A1 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A2 (.I(_0400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A3 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4242__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4223__A1 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4205__A2 (.I(_0403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A2 (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4207__I (.I(_0405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6541__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__A1 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__A2 (.I(_0406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4209__A2 (.I(_0407_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4241__A2 (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4218__I (.I(_0416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4344__A3 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4273__A2 (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4219__I (.I(_0417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4275__A2 (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4220__I (.I(_0418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7046__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__C1 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4229__A2 (.I(_0419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A3 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A1 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4228__A2 (.I(_0422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6821__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6820__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6815__A1 (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4225__I (.I(_0423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6786__A1 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A2 (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4226__I (.I(_0424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A2 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5121__I (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4862__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4227__A1 (.I(_0425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7072__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4448__A1 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4238__A2 (.I(_0434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4431__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4376__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4313__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A2 (.I(_0435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6509__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4339__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4268__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A1 (.I(_0438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4267__A2 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A3 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4244__A1 (.I(_0439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__B (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4259__A1 (.I(_0444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__A1 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4248__A2 (.I(_0445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4261__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4251__I (.I(_0448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A4 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4252__A2 (.I(_0449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A2 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__A3 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4254__C (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4253__A3 (.I(_0450_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A1 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4258__A2 (.I(_0455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I0 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A1 (.I(_0458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A3 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4341__A3 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4319__A2 (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4262__I (.I(_0459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4318__A2 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4282__A1 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4265__I (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4263__A3 (.I(_0460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4889__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A1 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4352__I (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4266__A3 (.I(_0463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__B1 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A2 (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4269__I (.I(_0466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A1 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4312__A2 (.I(_0467_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4271__A1 (.I(_0468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4306__B1 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4276__A2 (.I(_0469_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4305__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4274__A2 (.I(_0471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A2 (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4277__I (.I(_0474_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4880__A1 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4310__A2 (.I(_0475_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4877__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__A1 (.I(_0476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__B1 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4281__A2 (.I(_0477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A1 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4287__A2 (.I(_0480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__B1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6141__A1 (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4985__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4284__I (.I(_0481_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A1 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6167__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A2 (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4285__I (.I(_0482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6817__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5122__I (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4874__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4286__A1 (.I(_0483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A2 (.I(_0486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A1 (.I(_0487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4315__A4 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4297__A4 (.I(_0494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4346__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4345__A2 (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4298__I (.I(_0495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4872__I (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4300__A2 (.I(_0497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7042__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A1 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4303__A2 (.I(_0500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6823__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A1 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4308__A2 (.I(_0505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4311__A2 (.I(_0508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7074__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4450__A1 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4314__A2 (.I(_0510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A2 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A1 (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4317__I (.I(_0513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A1 (.I(_0515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4393__A3 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4320__A2 (.I(_0516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7115__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7114__B2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4324__A2 (.I(_0520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A1 (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4326__B (.I(_0522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4327__A2 (.I(_0523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4384__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4369__I (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4342__B (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A2 (.I(_0525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4332__B1 (.I(_0528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5701__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4385__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4336__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4335__A1 (.I(_0531_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A1 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4375__A2 (.I(_0537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__B1 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__A2 (.I(_0540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A2 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4348__B1 (.I(_0542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4410__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A3 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4355__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4347__A2 (.I(_0543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6873__A2 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A2 (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4349__I (.I(_0545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6571__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__A1 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4368__A2 (.I(_0546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5697__I (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I0 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4890__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4351__A1 (.I(_0547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__B1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B1 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4366__A2 (.I(_0549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A1 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4365__A2 (.I(_0550_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A3 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4402__A1 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A2 (.I(_0553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A1 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4364__A2 (.I(_0556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A2 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6175__A1 (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4362__I (.I(_0558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5123__I (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4363__A1 (.I(_0559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__B1 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5113__A3 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4408__I (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4371__A2 (.I(_0566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6867__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A2 (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4372__I (.I(_0568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6868__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6572__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A1 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4373__A2 (.I(_0569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7076__A1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4452__A1 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4377__A2 (.I(_0572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6577__I (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A2 (.I(_0574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5706__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A1 (.I(_0576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5076__A2 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4394__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4388__A1 (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4383__I (.I(_0578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A1 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A2 (.I(_0579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7119__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7116__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4386__A2 (.I(_0581_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__A2 (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4387__B (.I(_0582_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A1 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4430__A2 (.I(_0597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5135__A1 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A2 (.I(_0598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__B1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__B1 (.I(_0599_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4405__A2 (.I(_0600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A2 (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4407__I (.I(_0602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6585__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4906__A1 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4424__A2 (.I(_0603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7049__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4420__A2 (.I(_0604_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5590__A3 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__A1 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4412__A2 (.I(_0607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A1 (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5156__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4414__I (.I(_0609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6901__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A1 (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4415__I (.I(_0610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5195__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A2 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5118__I (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4416__A1 (.I(_0611_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A2 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5115__B (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4418__B1 (.I(_0613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4904__A1 (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4422__I (.I(_0617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7053__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4423__A1 (.I(_0618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4429__A2 (.I(_0620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6909__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6907__A2 (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4427__I (.I(_0622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6586__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4908__A1 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4428__A2 (.I(_0623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7078__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4454__A1 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4432__A2 (.I(_0626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4445__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4434__I (.I(_0628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4444__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4442__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A2 (.I(_0629_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4446__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4436__I (.I(_0630_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4443__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4441__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4439__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4437__A2 (.I(_0631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A1 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5923__A2 (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4456__I (.I(_0642_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A2 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5878__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A1 (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4457__I (.I(_0643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__B2 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A1 (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4459__I (.I(_0645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A1 (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4700__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4460__I (.I(_0646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5949__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A2 (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4462__I (.I(_0648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A2 (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5910__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4463__I (.I(_0649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__C2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A2 (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4464__I (.I(_0650_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4583__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A1 (.I(_0652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__B (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A1 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A2 (.I(_0653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__C (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A3 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A2 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A1 (.I(_0654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A1 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A2 (.I(_0655_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A2 (.I(_0656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__C (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4479__A2 (.I(_0657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__B2 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A1 (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4472__I (.I(_0658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5510__I (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A1 (.I(_0659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5441__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5437__I (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A1 (.I(_0660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A1 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4496__I (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A3 (.I(_0661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A1 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4476__A2 (.I(_0662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5780__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5014__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A2 (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4477__I (.I(_0663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5874__I (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4478__A2 (.I(_0664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A1 (.I(_0666_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A2 (.I(_0667_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5376__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5371__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A1 (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4482__I (.I(_0668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5029__I (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A1 (.I(_0669_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A2 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5454__I (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A1 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A3 (.I(_0670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A2 (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4485__I (.I(_0671_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5373__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A3 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A2 (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4486__I (.I(_0672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A1 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A3 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A3 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4487__A2 (.I(_0673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5802__A1 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A2 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__A3 (.I(_0674_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5213__I (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A1 (.I(_0675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5017__I (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4922__A2 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A1 (.I(_0676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A1 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4945__I (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4921__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4491__A2 (.I(_0677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A3 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A1 (.I(_0678_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5472__I (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A3 (.I(_0679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5473__I (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4494__A2 (.I(_0680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5457__A2 (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5367__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4495__I (.I(_0681_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__C (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A4 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5609__I (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B1 (.I(_0682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A1 (.I(_0683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5440__A2 (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4498__I (.I(_0684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__A2 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A3 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A3 (.I(_0685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6268__A1 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A2 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4501__B3 (.I(_0687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4582__A2 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4502__A3 (.I(_0688_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4559__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4530__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4506__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4504__I (.I(_0690_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4558__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__S (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4529__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4505__I (.I(_0691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4508__A2 (.I(_0692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A1 (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4707__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4511__I (.I(_0696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4513__A1 (.I(_0697_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A1 (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5970__B (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4515__I (.I(_0699_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A1 (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4516__I (.I(_0700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A1 (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4667__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4517__I (.I(_0701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4519__A1 (.I(_0702_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A2 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6028__A1 (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4521__I (.I(_0704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A1 (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4670__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4522__I (.I(_0705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4524__A1 (.I(_0706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6090__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6079__A1 (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4527__I (.I(_0709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6810__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A1 (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4673__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4528__I (.I(_0710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4637__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4599__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A1 (.I(_0711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4532__A2 (.I(_0712_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4542__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A2 (.I(_0713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6130__A1 (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4678__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4536__I (.I(_0717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4639__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4601__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4538__A1 (.I(_0718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6212__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6209__A1 (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6160__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4540__I (.I(_0720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A1 (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4681__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4541__I (.I(_0721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4641__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4603__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4543__A1 (.I(_0722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6220__A1 (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4722__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4546__I (.I(_0725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4685__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4643__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4605__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4548__A1 (.I(_0726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6272__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6253__A1 (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4551__I (.I(_0729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A1 (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4725__I (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4552__I (.I(_0730_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I0 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__I0 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__I0 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4553__I0 (.I(_0731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6343__A1 (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4688__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4557__I (.I(_0734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4649__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4611__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4561__A1 (.I(_0735_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6344__A1 (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4693__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4564__I (.I(_0740_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4651__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4613__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4566__A1 (.I(_0741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6415__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6372__A1 (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4568__I (.I(_0743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6367__A1 (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4734__I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4569__I (.I(_0744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4653__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4615__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4571__A1 (.I(_0745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A1 (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4737__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4574__I (.I(_0748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4655__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4617__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4576__A1 (.I(_0749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5400__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__A1 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4619__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A2 (.I(_0751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6107__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5905__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4579__I (.I(_0752_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__B1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__C2 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6393__B1 (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4581__I (.I(_0754_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6596__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A3 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__A2 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4584__A1 (.I(_0755_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4609__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4597__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4587__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4585__I (.I(_0758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4608__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4606__S (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4596__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4586__I (.I(_0759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4595__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4593__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4591__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4589__A2 (.I(_0760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4594__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4592__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4590__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4588__A2 (.I(_0761_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A2 (.I(_0774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6066__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6060__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5952__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4620__I (.I(_0780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__B1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__B1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__B1 (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4621__I (.I(_0781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5248__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4622__A2 (.I(_0782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4647__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4635__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4625__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4623__I (.I(_0783_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4646__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4644__S (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4634__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4624__I (.I(_0784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4633__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4631__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4629__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4627__A2 (.I(_0785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4632__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4626__A2 (.I(_0786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A2 (.I(_0799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__B1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__B1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__B1 (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4658__I (.I(_0805_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5904__B1 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5319__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4659__A2 (.I(_0806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4690__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4675__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4662__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4660__I (.I(_0807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4672__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4666__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4664__A2 (.I(_0809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4671__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4668__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4665__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4663__A2 (.I(_0810_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4669__A1 (.I(_0813_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5334__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5263__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4717__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4677__A1 (.I(_0817_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4684__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A2 (.I(_0819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5336__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5265__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4719__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4680__A1 (.I(_0821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5338__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5267__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4721__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4683__A1 (.I(_0823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4731__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A1 (.I(_0827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4699__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4697__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4692__A2 (.I(_0828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4733__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4695__A1 (.I(_0831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A1 (.I(_0835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4729__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4715__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4704__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4702__I (.I(_0836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4728__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__S (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4714__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4703__I (.I(_0837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4713__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4711__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4706__A2 (.I(_0838_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4712__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4710__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4708__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4705__A2 (.I(_0839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4709__A1 (.I(_0841_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4723__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4718__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4716__A2 (.I(_0846_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5340__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5269__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4724__A1 (.I(_0850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4736__A1 (.I(_0858_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4739__A1 (.I(_0860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5644__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__B (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A1 (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4741__I (.I(_0862_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A1 (.I(_0864_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4824__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4788__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4745__I (.I(_0866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A1 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4747__A2 (.I(_0868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__B (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5055__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A1 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A2 (.I(_0869_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A4 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A3 (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4749__I (.I(_0870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4795__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A2 (.I(_0871_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4893__A2 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4851__A1 (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4786__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4751__I (.I(_0872_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A4 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A2 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4772__I (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A3 (.I(_0875_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4816__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4755__I (.I(_0876_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4849__C (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4827__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A1 (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4756__I (.I(_0877_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6650__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6646__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5124__I (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4769__A1 (.I(_0879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A2 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4759__A1 (.I(_0880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A2 (.I(_0881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A2 (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4761__I (.I(_0882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5151__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5119__I (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5056__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A2 (.I(_0884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5020__I (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A3 (.I(_0885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4873__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A2 (.I(_0886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__B (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4766__I (.I(_0887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4887__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A2 (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__B (.I(_0889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A2 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4832__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__A1 (.I(_0892_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5097__I (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4953__I (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A1 (.I(_0893_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__B2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A2 (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4863__C (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__B (.I(_0895_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5522__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5146__I (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A1 (.I(_0896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__C (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A2 (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4776__C (.I(_0897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4828__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4814__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4808__I (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A2 (.I(_0900_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7107__A2 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A1 (.I(_0901_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A2 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4781__A1 (.I(_0902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4876__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A2 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__C (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__B1 (.I(_0903_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4879__A1 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4878__A2 (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__C (.I(_0904_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4784__B (.I(_0905_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__B (.I(_0911_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__I1 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__I1 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__I0 (.I(_0912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4792__A1 (.I(_0913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__B (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4809__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4793__I (.I(_0914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4902__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4901__B (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A2 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A1 (.I(_0915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4843__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4831__B (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4796__I (.I(_0917_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A2 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A1 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A4 (.I(_0920_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A1 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4909__A2 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4803__A3 (.I(_0921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A2 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4802__A4 (.I(_0923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4804__A2 (.I(_0925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__S (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4839__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4805__I (.I(_0926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A1 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4896__A2 (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__S (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4806__S (.I(_0927_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__B (.I(_0941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__I1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__I1 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I0 (.I(_0942_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4881__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__A2 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A1 (.I(_0944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4892__B (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4866__B (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4826__I (.I(_0945_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4837__A2 (.I(_0956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4838__B (.I(_0957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__S (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__S (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__S (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__S (.I(_0959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7112__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7105__A2 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A4 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__A1 (.I(_0961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4853__B (.I(_0971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4865__A1 (.I(_0975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7037__A2 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__B1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A4 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4864__A1 (.I(_0976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4886__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4861__A2 (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4860__I (.I(_0977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4869__B (.I(_0986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__I1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__I1 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4870__I0 (.I(_0987_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__B2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A2 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4903__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4875__A1 (.I(_0989_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4882__A2 (.I(_0997_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5430__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5296__A1 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4883__I0 (.I(_0999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4895__A2 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A1 (.I(_1001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4894__A2 (.I(_1008_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5298__I (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4897__A2 (.I(_1011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A2 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5508__I (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4900__A1 (.I(_1014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4910__A2 (.I(_1023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A1 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4911__I0 (.I(_1025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A1 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4914__A2 (.I(_1027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__C (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A2 (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4915__I (.I(_1028_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A1 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5792__I (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A2 (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4916__I (.I(_1029_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6071__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4927__A1 (.I(_1030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__B (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A2 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A3 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A1 (.I(_1031_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A1 (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5198__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4961__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4920__I (.I(_1033_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5036__I (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A1 (.I(_1034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A2 (.I(_1037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5377__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4925__A2 (.I(_1038_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A1 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4926__A2 (.I(_1039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7057__A2 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A1 (.I(_1042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A2 (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4931__I (.I(_1044_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5196__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4932__A2 (.I(_1045_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7102__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5194__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A1 (.I(_1046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5112__I (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A1 (.I(_1047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A1 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5105__I (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4935__A2 (.I(_1048_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A2 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4937__A1 (.I(_1050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5515__A1 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4938__A2 (.I(_1051_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5006__A1 (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__C (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4939__B (.I(_1052_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__A2 (.I(_1053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__C (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5442__A1 (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5372__I (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4941__I (.I(_1054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__B (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5871__I (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5065__A1 (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4942__I (.I(_1055_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6134__A1 (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4943__B (.I(_1056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A1 (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4946__I (.I(_1059_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A1 (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4947__I (.I(_1060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__B2 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5282__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A1 (.I(_1061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A3 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A4 (.I(_1062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5005__I (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A3 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A4 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A2 (.I(_1063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5854__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5847__A2 (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4951__I (.I(_1064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A2 (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__S (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4952__I (.I(_1065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A3 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4959__A2 (.I(_1066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__B (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4958__A1 (.I(_1067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A3 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4971__A2 (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4955__I (.I(_1068_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__A1 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5173__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A2 (.I(_1069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__A1 (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4957__I (.I(_1070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5519__A1 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A4 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4977__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A2 (.I(_1074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__B2 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A1 (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4962__I (.I(_1075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A1 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5535__I (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__C (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4963__A3 (.I(_1076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__C (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__B (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__C (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A1 (.I(_1078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5465__I (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5064__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4966__A2 (.I(_1079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5543__A2 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A1 (.I(_1080_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5565__B (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5381__I (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A1 (.I(_1081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A2 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A1 (.I(_1082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5558__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A1 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4970__A2 (.I(_1083_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A1 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5753__I (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A2 (.I(_1084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7141__A3 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A3 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A4 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4973__A3 (.I(_1086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__C (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7139__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4980__A2 (.I(_1087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5719__A2 (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5200__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4976__I (.I(_1089_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__B (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__C (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4979__A2 (.I(_1090_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A2 (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6500__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6453__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4978__I (.I(_1091_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__A1 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5000__A2 (.I(_1095_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5900__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A2 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4999__A1 (.I(_1096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5669__I (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__B (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__A1 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A2 (.I(_1097_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7085__A2 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__B (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4998__A1 (.I(_1098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6844__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6843__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6173__A1 (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4986__I (.I(_1099_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6850__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6849__A1 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__C2 (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4987__I (.I(_1100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6824__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__B1 (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4988__I (.I(_1101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A1 (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4989__I (.I(_1102_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A1 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__A2 (.I(_1103_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A1 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A2 (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4997__B (.I(_1105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5162__A4 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5050__A2 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A3 (.I(_1106_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5018__A2 (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4994__I (.I(_1107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7140__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A4 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A3 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4995__A2 (.I(_1108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7167__I (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7162__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4996__A2 (.I(_1109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7158__A1 (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__C (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__C (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5003__C (.I(_1116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__B2 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A1 (.I(_1117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6473__A4 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A1 (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5009__B (.I(_1121_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5030__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5019__I (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A1 (.I(_1123_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__B (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A1 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5012__A2 (.I(_1124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6655__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6449__I (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A1 (.I(_1125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6221__I (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5212__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A2 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A1 (.I(_1126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A1 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5015__A2 (.I(_1127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__B1 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5016__A2 (.I(_1128_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A3 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5024__A2 (.I(_1129_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5416__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A1 (.I(_1130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A2 (.I(_1131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A1 (.I(_1132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A1 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A2 (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5021__I (.I(_1133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A1 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5611__I (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5022__A2 (.I(_1134_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__B (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5023__A3 (.I(_1135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5661__A2 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A1 (.I(_1138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5846__A2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__A2 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5027__A3 (.I(_1139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A1 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5028__A2 (.I(_1140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__A2 (.I(_1141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A1 (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5031__I (.I(_1143_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A1 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5145__I (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A2 (.I(_1144_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__C (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__C (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A1 (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5033__I (.I(_1145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A1 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5040__I (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5034__A4 (.I(_1146_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5035__B1 (.I(_1147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5887__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5667__I (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A1 (.I(_1149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A3 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A3 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A3 (.I(_1150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6480__A3 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5899__I (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A1 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A4 (.I(_1151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__B (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A2 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__B1 (.I(_1152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A1 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__B2 (.I(_1153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5889__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5581__B (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A2 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A1 (.I(_1154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__A2 (.I(_1155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A2 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A3 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__B1 (.I(_1156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A1 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5363__I (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5045__B2 (.I(_1157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6468__C (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__C (.I(_1158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5069__A3 (.I(_1159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7117__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A2 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A1 (.I(_1160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5577__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5049__A1 (.I(_1161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A1 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5833__I (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5517__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__A2 (.I(_1162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A2 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5721__I (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B1 (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5051__B (.I(_1163_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A2 (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__C (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__B (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5059__B (.I(_1164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A2 (.I(_1166_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5058__A2 (.I(_1167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A3 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A3 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A1 (.I(_1168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__A2 (.I(_1169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6483__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A1 (.I(_1172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__B2 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5061__A1 (.I(_1173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A1 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5062__A2 (.I(_1174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A3 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5564__A1 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5063__A2 (.I(_1175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A3 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A2 (.I(_1176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5568__A2 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5068__A3 (.I(_1177_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7089__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__B1 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5066__A2 (.I(_1178_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__B1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5843__A1 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5067__A2 (.I(_1179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5205__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A1 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5141__A2 (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__B (.I(_1182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5144__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5085__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5072__A1 (.I(_1183_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5074__A4 (.I(_1186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__A2 (.I(_1187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__A2 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5079__A3 (.I(_1189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5082__B (.I(_1193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5084__A2 (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5083__C (.I(_1195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__B2 (.I(_1199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__B (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5088__I (.I(_1200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__A1 (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6540__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6512__I (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5089__C (.I(_1201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A1 (.I(_1202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5627__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A1 (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5091__I (.I(_1203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__C (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5713__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5597__A1 (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5092__I (.I(_1204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__B2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__B2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__B2 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5139__A1 (.I(_1205_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__A2 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5096__I1 (.I(_1208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__B (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__C (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__C (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5104__A2 (.I(_1210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6333__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6297__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A2 (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5099__I (.I(_1211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A2 (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5168__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5160__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5100__I (.I(_1212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5241__I (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B1 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5103__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5102__A2 (.I(_1214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__B (.I(_1217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6563__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6452__I (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5108__A1 (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5106__C (.I(_1218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__B2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__B2 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5109__A1 (.I(_1220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__A2 (.I(_1222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__B2 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__A1 (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5111__B (.I(_1223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5117__A2 (.I(_1228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5132__A2 (.I(_1230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6877__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6871__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A1 (.I(_1231_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__B (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__C (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5120__A2 (.I(_1232_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7083__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A1 (.I(_1234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A1 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A2 (.I(_1235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__B2 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A1 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5131__A3 (.I(_1236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A1 (.I(_1237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6691__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6682__A1 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5223__I (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A2 (.I(_1238_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A1 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5974__A2 (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5127__I (.I(_1239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6001__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5988__A1 (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5128__I (.I(_1240_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A1 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A3 (.I(_1241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A1 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5681__I (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5130__A4 (.I(_1242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5134__A2 (.I(_1246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A1 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5154__I (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5137__A2 (.I(_1249_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A2 (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5828__I (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5138__C (.I(_1250_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5140__A2 (.I(_1252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5193__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__A1 (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5143__I (.I(_1254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5203__A1 (.I(_1256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__C (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__C (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5528__I (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5149__A1 (.I(_1257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__C (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5726__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__A1 (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5147__I (.I(_1258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5703__I (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A2 (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5148__B (.I(_1259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__C (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6451__I (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5153__C (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5152__I (.I(_1263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__B (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__B (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__A2 (.I(_1264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__B1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5202__B1 (.I(_1265_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5676__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5655__I (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A2 (.I(_1266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__A2 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__B (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__A1 (.I(_1267_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6903__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A2 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A1 (.I(_1268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6814__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A1 (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5158__I (.I(_1269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6790__A1 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5177__I (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__B2 (.I(_1270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A1 (.I(_1271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6874__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6852__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6846__A1 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5164__B2 (.I(_1272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__C (.I(_1274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5175__A2 (.I(_1276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__B (.I(_1278_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6501__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A1 (.I(_1279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6299__A2 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6230__A1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__B1 (.I(_1280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__C (.I(_1282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__A2 (.I(_1283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5378__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5189__A2 (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5174__B (.I(_1284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A1 (.I(_1288_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A1 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A1 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5686__I (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__A2 (.I(_1289_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A1 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5182__B2 (.I(_1290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5491__A1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__B1 (.I(_1292_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6590__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__A1 (.I(_1295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6562__A1 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5188__B2 (.I(_1296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6758__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5495__I (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__B1 (.I(_1298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7138__A1 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A3 (.I(_1301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A1 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5245__I (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5197__A2 (.I(_1307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A1 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__B2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__B2 (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5199__B (.I(_1310_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__B (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__C (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__C (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5201__B (.I(_1312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5204__A2 (.I(_1315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A2 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5211__I (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A1 (.I(_1317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__C (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A2 (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5208__I (.I(_1318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7079__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5209__A2 (.I(_1319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A2 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A1 (.I(_1321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__A1 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A3 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A2 (.I(_1322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A1 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5218__A3 (.I(_1323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5992__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5879__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5370__I (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5214__A1 (.I(_1324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5894__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5785__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__A2 (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5215__I (.I(_1325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__C (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A1 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5922__A2 (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5216__I (.I(_1326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A1 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5982__I (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__B (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5217__A2 (.I(_1327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5225__A2 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5220__I (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5219__A1 (.I(_1329_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5221__A2 (.I(_1331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5224__A1 (.I(_1333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5358__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5233__A1 (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5228__I (.I(_1336_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5990__I (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A1 (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5229__I (.I(_1337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5888__A2 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5232__A1 (.I(_1338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5239__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5231__A2 (.I(_1339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A3 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5606__A3 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A3 (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5234__I (.I(_1341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5459__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5380__A2 (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5235__I (.I(_1342_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5945__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A3 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5364__A2 (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5236__I (.I(_1343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__A2 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A1 (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5237__I (.I(_1344_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__A2 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__B1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5238__A1 (.I(_1345_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5240__A2 (.I(_1346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6853__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6847__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A1 (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5242__I (.I(_1348_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5243__A1 (.I(_1349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5841__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5840__A2 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5246__A1 (.I(_1351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5273__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5261__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5251__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5249__I (.I(_1353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5272__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5270__S (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5260__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5250__I (.I(_1354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5259__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5257__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5255__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5253__A2 (.I(_1355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5258__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5256__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A2 (.I(_1356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A2 (.I(_1362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5281__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5279__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5277__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5275__A2 (.I(_1368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5288__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5283__I (.I(_1374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5301__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5299__A2 (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5286__S (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5284__S (.I(_1375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5295__I (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5293__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__S (.I(_1378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5344__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5332__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5322__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5320__I (.I(_1395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5343__I (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5341__S (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5331__I (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5321__I (.I(_1396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5330__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5328__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5326__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5324__A2 (.I(_1397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5327__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A2 (.I(_1398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5352__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5350__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5348__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5346__A2 (.I(_1410_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6223__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A2 (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5366__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5354__I (.I(_1416_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5626__A1 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A2 (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5355__I (.I(_1417_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6860__A2 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A1 (.I(_1418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5447__A1 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A2 (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5357__I (.I(_1419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__B2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A1 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A2 (.I(_1420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__B (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5359__I (.I(_1421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__B (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A3 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5857__A3 (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5360__I (.I(_1422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6037__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A2 (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5776__I (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5361__I (.I(_1423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__B2 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__B (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5362__A3 (.I(_1424_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A2 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A1 (.I(_1426_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__B (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__B2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5365__A2 (.I(_1427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6892__I (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__B2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__B2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__A2 (.I(_1428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6799__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__A2 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A1 (.I(_1429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6002__A2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__B2 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A3 (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5368__I (.I(_1430_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5882__A1 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5598__I (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__A2 (.I(_1431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A1 (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5375__B (.I(_1432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A1 (.I(_1433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6737__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__A1 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A2 (.I(_1434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__C (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__C (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__C (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A3 (.I(_1435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A1 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A3 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5374__A4 (.I(_1436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5978__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5714__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5403__I (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5383__A1 (.I(_1439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5562__B (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A1 (.I(_1440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A2 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5379__A2 (.I(_1441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A1 (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5534__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5524__I (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5382__C (.I(_1444_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5384__A2 (.I(_1446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5521__A1 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5386__A2 (.I(_1448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5480__I (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A2 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5387__A4 (.I(_1449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5640__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5389__A1 (.I(_1451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6040__I (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5391__A2 (.I(_1453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A1 (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6072__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5545__I (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5393__B (.I(_1455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A2 (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5394__C (.I(_1456_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A2 (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5395__I (.I(_1457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6896__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6710__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5407__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5397__I (.I(_1459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__B (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5707__I (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5398__I (.I(_1460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__B (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__B (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__B (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5399__B (.I(_1461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__C (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__B (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__B (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5402__B (.I(_1463_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__C (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__C (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__A1 (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5404__I (.I(_1465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7080__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6559__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5794__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5405__A1 (.I(_1466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5817__B (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__B (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5414__B (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__B (.I(_1470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6430__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5912__A1 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5413__A2 (.I(_1473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5422__I (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5417__I (.I(_1476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5434__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5432__A2 (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5420__S (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5418__S (.I(_1477_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5429__I (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5427__S (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5425__S (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5423__S (.I(_1480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5488__A1 (.I(_1488_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5718__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5624__I (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5438__A1 (.I(_1489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5762__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5439__A2 (.I(_1490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5630__A2 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A1 (.I(_1491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5789__I (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A1 (.I(_1494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5452__A2 (.I(_1499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6732__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6442__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5735__I (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5451__A1 (.I(_1500_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A1 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6675__I (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5450__A2 (.I(_1501_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5453__A2 (.I(_1504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A1 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5462__I (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5456__A2 (.I(_1506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6630__A1 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A2 (.I(_1508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__C (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5458__A2 (.I(_1509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6660__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5893__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5749__I (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5470__A2 (.I(_1511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6137__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A2 (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5461__I (.I(_1512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__A2 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A1 (.I(_1513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A1 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5752__I (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5463__A2 (.I(_1514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__C (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B1 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5541__I (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A2 (.I(_1516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5850__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A1 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5623__A2 (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5466__I (.I(_1517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__B2 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5549__A2 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5542__B2 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A3 (.I(_1518_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__B (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6556__A1 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5646__I (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A2 (.I(_1519_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__B1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__B1 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A4 (.I(_1520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5853__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__A1 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A2 (.I(_1523_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5566__A2 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A1 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A3 (.I(_1524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6049__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5983__I (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A3 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A4 (.I(_1525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A1 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A2 (.I(_1526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5576__A1 (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5476__I (.I(_1527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5642__A2 (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5478__I (.I(_1529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A2 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5759__I (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A3 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5479__A2 (.I(_1530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5574__B (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5482__A4 (.I(_1533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5483__A4 (.I(_1534_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5501__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5499__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5486__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5484__I (.I(_1535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6912__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6906__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5487__A1 (.I(_1537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__A2 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6932__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6306__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5490__A1 (.I(_1540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6342__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5493__A1 (.I(_1542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7081__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5498__A1 (.I(_1544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A2 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5497__A1 (.I(_1545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5507__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5505__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5503__A2 (.I(_1547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6404__A3 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A1 (.I(_1548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5502__A2 (.I(_1549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6876__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6870__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A1 (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5509__I (.I(_1553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__B2 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5512__A1 (.I(_1554_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5625__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5575__B2 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5511__A1 (.I(_1555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5546__A2 (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5514__I (.I(_1557_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6631__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6467__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5569__A1 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A2 (.I(_1558_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5516__A4 (.I(_1559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6178__I (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A2 (.I(_1562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5594__I (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5520__A3 (.I(_1563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__B2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5527__A2 (.I(_1564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7091__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A1 (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5523__I (.I(_1566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5693__A2 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__A1 (.I(_1567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5711__I (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5643__A1 (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5525__C (.I(_1568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5526__A2 (.I(_1569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__A1 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A2 (.I(_1571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7131__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__C (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5529__A1 (.I(_1572_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__C (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__C (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__C (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5533__C (.I(_1576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__C (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5747__I (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5544__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A1 (.I(_1577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__A1 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5699__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A2 (.I(_1578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7090__A1 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__A2 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5537__A3 (.I(_1579_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__B (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__B (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__B2 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__A1 (.I(_1583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5582__A1 (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5552__B (.I(_1584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A1 (.I(_1585_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A1 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5551__A2 (.I(_1586_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__C (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__C (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__C (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A1 (.I(_1587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6672__I (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5773__A2 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A4 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5548__A2 (.I(_1589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A2 (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__B (.I(_1590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__C (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5641__A2 (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5550__C (.I(_1591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5555__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A2 (.I(_1594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__C (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__C (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5746__I (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__B (.I(_1595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5716__I (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5559__A1 (.I(_1598_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5851__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5560__A2 (.I(_1600_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5561__A2 (.I(_1601_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6636__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A1 (.I(_1602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5724__I (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5563__A2 (.I(_1603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5586__A2 (.I(_1605_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5849__A1 (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5567__C (.I(_1607_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A1 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__B (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A2 (.I(_1609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5845__A2 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5570__A3 (.I(_1610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6632__A3 (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5572__I (.I(_1612_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5865__A2 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5651__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5593__I (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5573__A4 (.I(_1613_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A1 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A2 (.I(_1615_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A2 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6653__I (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A1 (.I(_1617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6465__B1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A1 (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5578__I (.I(_1618_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__B (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__B (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__B2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__A2 (.I(_1619_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7014__B (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A2 (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__B (.I(_1620_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A1 (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5583__C (.I(_1623_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5584__A4 (.I(_1624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5585__A2 (.I(_1625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A1 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A2 (.I(_1628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5748__A3 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5725__A2 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5591__A4 (.I(_1631_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6637__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5622__A1 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5592__A2 (.I(_1632_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5605__A1 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A2 (.I(_1633_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__B2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A2 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5603__A1 (.I(_1634_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A3 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5602__A2 (.I(_1635_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5739__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A2 (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5596__I (.I(_1636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5808__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__B (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A1 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A2 (.I(_1637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__C (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5599__A1 (.I(_1639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__B2 (.I(_1640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5698__I (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A2 (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__C (.I(_1641_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A2 (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5608__C (.I(_1647_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5859__A1 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5616__A2 (.I(_1648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A3 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5728__A1 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5610__A2 (.I(_1649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7159__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__A1 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A2 (.I(_1651_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A1 (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5613__I (.I(_1652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5614__A1 (.I(_1653_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A1 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5615__A4 (.I(_1654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A4 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5660__A2 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5618__A4 (.I(_1657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A1 (.I(_1658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5620__A2 (.I(_1659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A1 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5621__A4 (.I(_1660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A1 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A2 (.I(_1662_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5848__C (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A1 (.I(_1663_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A2 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5632__A1 (.I(_1664_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A2 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5723__C (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__B1 (.I(_1665_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5629__C (.I(_1668_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A2 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A4 (.I(_1670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5633__A2 (.I(_1672_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5635__A2 (.I(_1673_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A2 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__B (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A1 (.I(_1675_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6718__I (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5738__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5638__A2 (.I(_1676_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6826__B (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6765__I (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5639__A2 (.I(_1677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A2 (.I(_1682_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6888__I (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5645__A2 (.I(_1683_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5860__A1 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5648__A3 (.I(_1684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6527__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6446__I (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5647__A1 (.I(_1685_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A2 (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__B (.I(_1687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6863__B (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6829__A1 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A2 (.I(_1689_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7170__C (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__C (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__C (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__C (.I(_1691_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7153__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7122__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7097__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5657__A2 (.I(_1692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7103__A1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I1 (.I(_1694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A3 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5662__A2 (.I(_1698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5696__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A1 (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5664__I (.I(_1700_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__S (.I(_1701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5668__A2 (.I(_1703_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A1 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5689__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5683__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A2 (.I(_1705_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__B (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7157__A1 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5671__A2 (.I(_1706_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I1 (.I(_1707_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__A2 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A1 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5679__A2 (.I(_1709_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7034__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5678__A1 (.I(_1710_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A1 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A2 (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5677__I (.I(_1711_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__B2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5680__A2 (.I(_1713_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7147__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5682__A1 (.I(_1715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A2 (.I(_1716_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__B (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7151__A1 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5684__A3 (.I(_1717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5685__B (.I(_1718_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6788__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__A1 (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5687__I (.I(_1719_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7137__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5688__A1 (.I(_1720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__B (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7145__A1 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5690__A2 (.I(_1722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5691__I1 (.I(_1723_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A2 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5694__I1 (.I(_1725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7050__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A1 (.I(_1728_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7176__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7163__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__A1 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5700__A2 (.I(_1729_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5702__A2 (.I(_1731_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A1 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5704__A2 (.I(_1733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5705__A2 (.I(_1734_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7126__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__B (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__B (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5709__A1 (.I(_1736_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5830__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5712__A1 (.I(_1739_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7082__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6566__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A1 (.I(_1741_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5730__A1 (.I(_1743_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7087__A2 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6439__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6341__A3 (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5717__I (.I(_1744_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__A2 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__A1 (.I(_1745_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5727__A2 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A3 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B1 (.I(_1746_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5764__A2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5720__B2 (.I(_1747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__C (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6198__I (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__C (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5722__A2 (.I(_1749_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5729__A1 (.I(_1751_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5731__B1 (.I(_1758_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5732__A2 (.I(_1759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5743__A2 (.I(_1760_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6795__C (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6513__I (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5740__B (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5736__I (.I(_1763_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A1 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A2 (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5737__B (.I(_1764_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5742__B1 (.I(_1765_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A3 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5741__A4 (.I(_1768_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__A2 (.I(_1771_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7136__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7101__B (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6746__A1 (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5745__B (.I(_1772_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6293__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6251__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5821__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A1 (.I(_1773_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__C (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__C (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5771__I (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A1 (.I(_1774_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__B2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A1 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5869__B (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__A2 (.I(_1775_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__B2 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5811__A3 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5750__A1 (.I(_1776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__B1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5761__A1 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5757__B2 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A4 (.I(_1778_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__A2 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A2 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5812__I (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A1 (.I(_1779_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__B2 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A1 (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5754__I (.I(_1780_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5765__B2 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5755__A1 (.I(_1781_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5756__A2 (.I(_1782_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A2 (.I(_1784_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__C (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__C (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A1 (.I(_1785_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A1 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6883__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__B2 (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5760__I (.I(_1786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__B (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__C (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__C (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5763__A1 (.I(_1787_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__A3 (.I(_1790_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5767__B (.I(_1793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5768__A3 (.I(_1794_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5769__B (.I(_1795_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5770__A2 (.I(_1796_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__A2 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__A1 (.I(_1797_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__C (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__B (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__C (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__B (.I(_1798_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6208__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6171__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5980__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5774__I (.I(_1799_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6436__B (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6400__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5915__B (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A1 (.I(_1801_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6383__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__B2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__B2 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A1 (.I(_1802_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5788__B (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5784__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A2 (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__B (.I(_1803_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5779__A3 (.I(_1804_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6269__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6222__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6099__A2 (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5781__I (.I(_1806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A2 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6235__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5782__A1 (.I(_1807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__B (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5783__A2 (.I(_1808_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__A2 (.I(_1809_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__A2 (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6048__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5786__I (.I(_1811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6352__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A1 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5787__B2 (.I(_1812_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__B1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__B1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5790__A1 (.I(_1815_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A1 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A2 (.I(_1818_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__A2 (.I(_1820_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5796__B1 (.I(_1821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5797__C (.I(_1822_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5816__A2 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5800__A1 (.I(_1823_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5805__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5801__A2 (.I(_1825_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__B1 (.I(_1827_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__C (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__C (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__B1 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A2 (.I(_1828_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__C (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6696__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5825__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5807__I (.I(_1831_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__A1 (.I(_1832_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__B (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__B2 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6505__A1 (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5810__B (.I(_1834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__B1 (.I(_1836_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6545__A2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5813__B2 (.I(_1837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5824__A2 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5823__A3 (.I(_1844_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__C (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__A1 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5835__A3 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A3 (.I(_1847_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6667__A1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__B1 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5829__A2 (.I(_1850_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5844__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5832__C (.I(_1853_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6546__A2 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__B1 (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5834__I (.I(_1854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__B1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6582__B1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__A2 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5837__A1 (.I(_1855_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6635__A3 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A2 (.I(_1868_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5852__B (.I(_1870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6455__I (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5855__A2 (.I(_1873_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6634__A4 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5856__A3 (.I(_1874_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__B (.I(_1879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5862__A4 (.I(_1880_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5867__I (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5863__I (.I(_1881_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6116__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5968__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5917__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5864__I (.I(_1882_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6438__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6402__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5916__A2 (.I(_1883_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5921__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5866__I (.I(_1884_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A1 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__A2 (.I(_1885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__C (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__C (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__C (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5868__B (.I(_1886_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6163__I (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5870__I (.I(_1888_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6424__A1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__A1 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5972__I (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__A2 (.I(_1889_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6349__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6183__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5876__A1 (.I(_1890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6273__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5873__A1 (.I(_1891_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__B2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A1 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__A2 (.I(_1896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__B2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__B2 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A1 (.I(_1897_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A1 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5880__A2 (.I(_1898_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A2 (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5881__B (.I(_1899_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5885__A2 (.I(_1902_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5892__B (.I(_1906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6218__I (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6050__I (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__B2 (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5890__I (.I(_1908_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A1 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A1 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5995__A1 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5891__A4 (.I(_1909_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5898__B1 (.I(_1912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A1 (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5895__I (.I(_1913_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A1 (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6086__I (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5896__I (.I(_1914_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A1 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__B2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__B2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5897__A2 (.I(_1915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7012__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__A1 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6247__B (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__A2 (.I(_1918_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__B2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__B2 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5913__A1 (.I(_1919_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6283__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6109__A1 (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__B (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5903__I (.I(_1921_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6433__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6245__B2 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5962__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5908__A1 (.I(_1922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A2 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__B1 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__A2 (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5906__I (.I(_1924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__B1 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5907__B2 (.I(_1925_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6429__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A2 (.I(_1929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5914__B (.I(_1932_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6364__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6329__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6206__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5966__A2 (.I(_1936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A2 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5920__A1 (.I(_1937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5965__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__A2 (.I(_1938_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__B2 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__C (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5964__A1 (.I(_1939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6080__I (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5973__I (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A1 (.I(_1940_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5947__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5936__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5932__A2 (.I(_1941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6703__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5934__A1 (.I(_1944_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5931__A2 (.I(_1948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5933__A2 (.I(_1950_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5935__C (.I(_1952_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A2 (.I(_1956_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A1 (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5942__B (.I(_1959_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5943__B2 (.I(_1960_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5944__A3 (.I(_1961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5946__A1 (.I(_1963_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A1 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__C (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__C (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__B2 (.I(_1966_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__A2 (.I(_1968_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__A2 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__B1 (.I(_1969_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6240__I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6008__I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5957__I (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__A2 (.I(_1970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6241__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6010__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5958__I (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5954__B1 (.I(_1971_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__B1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__B1 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A2 (.I(_1975_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__B1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__B1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__B1 (.I(_1976_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__A2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__B1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__B1 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__C2 (.I(_1977_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5963__C (.I(_1980_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6159__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6115__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6077__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6024__A2 (.I(_1984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6292__A2 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__A1 (.I(_1985_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6117__A3 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6078__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A2 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5971__A1 (.I(_1986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__A1 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__A2 (.I(_1988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A2 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__B1 (.I(_1994_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__C (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__C (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__C (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5979__C (.I(_1995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6923__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__A1 (.I(_2000_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5985__A2 (.I(_2001_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6954__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6345__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5989__A1 (.I(_2003_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5994__A2 (.I(_2006_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5991__A1 (.I(_2007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5993__A1 (.I(_2009_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__A2 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A1 (.I(_2013_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6042__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6041__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6000__A2 (.I(_2014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__A2 (.I(_2017_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6405__C (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__B (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__C (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6004__C (.I(_2020_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6005__B (.I(_2021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6006__A2 (.I(_2022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6019__A2 (.I(_2023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6149__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6105__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6065__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6012__A1 (.I(_2024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6015__A2 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6009__B1 (.I(_2025_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__B1 (.I(_2027_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__B (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6153__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6070__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6016__A1 (.I(_2030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6018__B1 (.I(_2034_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__B2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__B2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__B2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6021__B2 (.I(_2037_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6114__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6076__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6023__B (.I(_2039_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6026__A1 (.I(_2041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6075__A1 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6053__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__A2 (.I(_2042_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6029__A1 (.I(_2043_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6054__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6034__A2 (.I(_2049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__B2 (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6035__B (.I(_2050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6236__C (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6038__I (.I(_2053_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A1 (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6039__B (.I(_2054_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A1 (.I(_2056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6096__A2 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6045__A2 (.I(_2060_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6047__A2 (.I(_2062_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__A2 (.I(_2063_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A1 (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6058__B (.I(_2064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6229__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__B2 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6057__A1 (.I(_2065_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__A1 (.I(_2066_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6089__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6052__A2 (.I(_2067_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6056__B2 (.I(_2071_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6074__A2 (.I(_2074_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__A2 (.I(_2075_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__B1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__A2 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B1 (.I(_2076_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__B1 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__A2 (.I(_2078_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__B1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__B1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__B1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6064__B1 (.I(_2079_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__B1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A2 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__B1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6067__B1 (.I(_2082_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__B1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__B1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__B1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6069__B1 (.I(_2084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__B (.I(_2087_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__C (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__B (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__C (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6073__C (.I(_2088_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6113__A1 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6091__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__A2 (.I(_2094_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6260__A3 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6084__A2 (.I(_2098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6801__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__A2 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B1 (.I(_2100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__B2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__B2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__B2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6087__B2 (.I(_2101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__A2 (.I(_2105_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__C (.I(_2107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6094__B1 (.I(_2108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6139__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6138__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A2 (.I(_2110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6140__A1 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6098__A3 (.I(_2112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__A2 (.I(_2113_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A2 (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6100__B (.I(_2114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6101__B (.I(_2115_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6102__A2 (.I(_2116_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6112__A2 (.I(_2117_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6284__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__B1 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A2 (.I(_2122_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6110__A3 (.I(_2124_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6111__B (.I(_2125_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6158__A1 (.I(_2130_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6157__A1 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6133__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__A2 (.I(_2132_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6129__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6123__A1 (.I(_2135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6132__A2 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6125__B1 (.I(_2138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6834__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6161__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A1 (.I(_2141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6219__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A2 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6131__A1 (.I(_2142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__A2 (.I(_2145_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6136__B2 (.I(_2149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A1 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__B (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__A2 (.I(_2151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6143__A2 (.I(_2156_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6144__C (.I(_2157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6145__B (.I(_2158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6156__A2 (.I(_2160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6354__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6318__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A2 (.I(_2164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6155__B1 (.I(_2168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6180__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6162__A1 (.I(_2173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__A1 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A2 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6182__A2 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__A2 (.I(_2175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6181__A2 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6170__B1 (.I(_2182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6231__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6177__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6176__A1 (.I(_2187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A1 (.I(_2190_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6966__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6830__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6769__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6179__A2 (.I(_2191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6186__A2 (.I(_2192_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6185__B2 (.I(_2197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6187__A2 (.I(_2199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__A1 (.I(_2201_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6285__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6282__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A2 (.I(_2206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6358__B (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6323__B (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6286__A1 (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6197__B (.I(_2209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__B (.I(_2210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6397__B (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__C (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B2 (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6199__C (.I(_2211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6200__B (.I(_2212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__B2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__B2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__B2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6203__B2 (.I(_2215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6363__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6328__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6205__B (.I(_2217_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6307__A2 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6271__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6250__A1 (.I(_2219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6925__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6833__C (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6249__A1 (.I(_2220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6248__I (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6225__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__A2 (.I(_2222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6215__A2 (.I(_2226_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__C (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6216__B (.I(_2227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A2 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6228__A1 (.I(_2230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6380__B (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__C (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__B (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A1 (.I(_2233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A2 (.I(_2234_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6891__A1 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6224__A3 (.I(_2235_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6234__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6233__A2 (.I(_2244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6237__A3 (.I(_2248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__B1 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__A2 (.I(_2252_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__B1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6428__B1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6392__B1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6244__B1 (.I(_2253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6246__B1 (.I(_2257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6291__B2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6276__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6264__A2 (.I(_2264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6275__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6263__A2 (.I(_2273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6267__B (.I(_2277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6279__A2 (.I(_2281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6278__A2 (.I(_2283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6922__A1 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6274__A2 (.I(_2284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6277__A2 (.I(_2285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6280__A2 (.I(_2290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6287__A2 (.I(_2294_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6288__B (.I(_2298_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6944__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6308__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6296__A1 (.I(_2304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6327__A1 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6310__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__A2 (.I(_2306_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6960__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6939__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6413__A2 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6302__A1 (.I(_2308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6309__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6303__A2 (.I(_2312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6943__A1 (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6304__B (.I(_2313_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6326__A1 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6305__A2 (.I(_2314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6316__A2 (.I(_2316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6315__A2 (.I(_2318_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6934__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A2 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6340__I (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6312__A1 (.I(_2321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__B (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6313__A2 (.I(_2322_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6314__B1 (.I(_2323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6317__A2 (.I(_2326_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6324__B (.I(_2333_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6325__B (.I(_2334_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6374__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6373__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6365__I (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6332__A1 (.I(_2339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6362__A1 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6348__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__A2 (.I(_2341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6347__A2 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6338__B1 (.I(_2346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6351__A2 (.I(_2351_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__A2 (.I(_2353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6346__A2 (.I(_2354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6350__B1 (.I(_2355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6359__B (.I(_2367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6360__B (.I(_2368_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A2 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6366__A1 (.I(_2373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__A2 (.I(_2375_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6388__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6378__A2 (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6370__I (.I(_2377_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6401__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__A2 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6371__B1 (.I(_2378_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6985__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6391__B1 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6379__A2 (.I(_2385_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6382__A4 (.I(_2389_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A1 (.I(_2392_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6403__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6387__A2 (.I(_2394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6389__A2 (.I(_2395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6390__A3 (.I(_2397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6394__A2 (.I(_2400_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6398__B2 (.I(_2405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6399__B (.I(_2406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6427__A1 (.I(_2412_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6410__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6407__A1 (.I(_2413_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6437__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6419__A2 (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6409__I (.I(_2415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6412__A3 (.I(_2418_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6425__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6420__A2 (.I(_2425_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7005__A1 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6422__A3 (.I(_2428_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6423__A4 (.I(_2429_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__C (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6426__C (.I(_2432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6434__A3 (.I(_2440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6435__B (.I(_2441_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6921__A1 (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6494__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6440__I (.I(_2445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6987__A2 (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6539__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__C (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6441__I (.I(_2446_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6854__C (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6764__C (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6692__C (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6443__I (.I(_2448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__B2 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A1 (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6444__I (.I(_2449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6487__A1 (.I(_2454_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__C (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6803__A1 (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__B (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__B (.I(_2455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6580__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6551__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6461__A2 (.I(_2457_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__B1 (.I(_2460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6547__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A2 (.I(_2461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7086__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6564__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6460__A1 (.I(_2465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A2 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6484__A1 (.I(_2468_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6818__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6756__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6678__I (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A2 (.I(_2476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6479__B (.I(_2479_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6475__A3 (.I(_2480_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6952__A1 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6949__B (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__C (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6477__A2 (.I(_2482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6482__A1 (.I(_2486_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6553__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6492__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6488__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6485__I (.I(_2490_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A1 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6537__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6524__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A2 (.I(_2494_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7188__B (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7152__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7146__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6508__A1 (.I(_2496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A1 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A2 (.I(_2497_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6557__C (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6528__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6497__A1 (.I(_2499_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6507__B1 (.I(_2502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B1 (.I(_2507_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6504__B2 (.I(_2508_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6506__A2 (.I(_2510_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__A2 (.I(_2515_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__C (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6558__B (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6529__B (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6516__B (.I(_2516_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__C (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__B2 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6526__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A1 (.I(_2517_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A2 (.I(_2520_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__B (.I(_2521_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__C (.I(_2522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6523__A3 (.I(_2525_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6525__A1 (.I(_2527_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6536__A2 (.I(_2532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7174__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6531__A1 (.I(_2533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6534__B1 (.I(_2535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__C (.I(_2537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6772__A1 (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6588__B (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6574__B (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6544__B (.I(_2542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__A1 (.I(_2546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6550__A2 (.I(_2551_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6552__A4 (.I(_2553_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6554__A2 (.I(_2555_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6555__B (.I(_2556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__B (.I(_2559_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7084__A1 (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6589__B (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6575__B (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__B (.I(_2561_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__B1 (.I(_2563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6565__B2 (.I(_2565_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6567__C (.I(_2567_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__A2 (.I(_2568_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__B (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6594__B (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6583__B (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6569__B (.I(_2569_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6570__B (.I(_2570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6584__A1 (.I(_2574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A1 (.I(_2576_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__B1 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7054__A2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6593__B2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6578__A2 (.I(_2577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6579__A2 (.I(_2578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6581__A2 (.I(_2580_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6591__B2 (.I(_2589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6592__A2 (.I(_2590_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6595__A2 (.I(_2592_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6621__I (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6609__I (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6599__I (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6597__I (.I(_2594_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6620__I (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6618__S (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6608__I (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6598__I (.I(_2595_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6607__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6605__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6603__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6601__A2 (.I(_2596_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6606__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A2 (.I(_2597_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6617__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6615__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6613__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6611__A2 (.I(_2602_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6616__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6614__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6612__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6610__A2 (.I(_2603_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6629__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6627__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6625__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6623__A2 (.I(_2609_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6628__A2 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6626__A2 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6624__A2 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6622__A2 (.I(_2610_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A1 (.I(_2616_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6633__A2 (.I(_2617_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6743__I (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6638__I (.I(_2622_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A2 (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6640__I (.I(_2624_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6807__A1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6775__A1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6712__A1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6671__A1 (.I(_2625_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A1 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__B (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6677__A2 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A1 (.I(_2626_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6819__C (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6725__B (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6683__I (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6643__I (.I(_2627_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6935__A1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6913__B2 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__C (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6651__A1 (.I(_2628_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6657__A2 (.I(_2636_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A2 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6661__A1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A1 (.I(_2637_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A1 (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6654__I (.I(_2638_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A1 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__B2 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__A2 (.I(_2639_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__B (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__C (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__B (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6656__C (.I(_2640_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6663__B (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6659__I (.I(_2643_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__B2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__B2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__B2 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__A1 (.I(_2644_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__B1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__B1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6800__A1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__B1 (.I(_2645_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6662__B2 (.I(_2646_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6858__I (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__A2 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6700__I (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6664__B1 (.I(_2648_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6665__A2 (.I(_2649_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6894__A2 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6804__A2 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6668__B1 (.I(_2652_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6670__A2 (.I(_2654_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__B2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6708__I (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6673__A2 (.I(_2656_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6808__I (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__A2 (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6674__I (.I(_2657_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6864__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__A2 (.I(_2658_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A1 (.I(_2659_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6702__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6695__A2 (.I(_2660_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A1 (.I(_2661_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6904__A1 (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6762__B (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6730__B (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6687__I (.I(_2670_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6694__A2 (.I(_2677_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6707__A1 (.I(_2679_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6919__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6768__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6699__A1 (.I(_2680_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6968__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6771__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6706__A2 (.I(_2684_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6704__B2 (.I(_2687_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6970__B2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6926__B2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6773__B2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6709__B2 (.I(_2692_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__B (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__B (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6774__B (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__B (.I(_2694_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6992__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6972__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6836__A1 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A2 (.I(_2696_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6739__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6736__A2 (.I(_2698_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__B (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6981__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A1 (.I(_2701_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6784__B1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6754__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6724__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__A1 (.I(_2704_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__B (.I(_2714_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__B (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__B (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6825__C (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6733__C (.I(_2715_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6735__A2 (.I(_2717_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__B2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__B2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__B2 (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6738__B (.I(_2720_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6924__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6802__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6741__A2 (.I(_2721_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6740__B2 (.I(_2722_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6742__B1 (.I(_2724_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__B1 (.I(_2725_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7007__C (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6837__I (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6835__A2 (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6744__C (.I(_2726_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6770__A2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__A2 (.I(_2733_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6936__A1 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__B2 (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6855__B (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6766__B (.I(_2747_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6767__B (.I(_2748_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6777__A2 (.I(_2757_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__A2 (.I(_2759_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6798__A2 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__B1 (.I(_2762_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6787__A2 (.I(_2767_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A1 (.I(_2769_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6796__A2 (.I(_2776_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6797__C (.I(_2777_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6927__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6897__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6806__A2 (.I(_2786_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__A2 (.I(_2791_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6831__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__A2 (.I(_2793_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6827__B (.I(_2806_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6828__B (.I(_2807_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6832__B1 (.I(_2811_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6946__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6928__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6898__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6866__A1 (.I(_2816_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__A2 (.I(_2819_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6859__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__A2 (.I(_2821_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6856__B (.I(_2834_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6857__B (.I(_2835_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__A2 (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__A2 (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__A2 (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6862__A2 (.I(_2837_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6861__B2 (.I(_2839_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6872__A2 (.I(_2848_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6878__A2 (.I(_2854_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6885__A2 (.I(_2857_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6890__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6884__A2 (.I(_2860_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__B (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__B (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__B (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6889__B (.I(_2866_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__B2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__B2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6942__B2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6893__B2 (.I(_2870_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6947__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6933__A2 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6905__A1 (.I(_2879_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A2 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A1 (.I(_2885_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6951__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6948__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6931__A3 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6911__A2 (.I(_2887_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6914__B1 (.I(_2890_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6920__B (.I(_2896_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6941__A2 (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__A2 (.I(_2906_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6937__B (.I(_2912_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6940__A2 (.I(_2915_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A3 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__B (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A2 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A1 (.I(_2922_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__C (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A2 (.I(_2923_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6950__A3 (.I(_2924_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6975__A2 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6953__A1 (.I(_2926_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6958__A2 (.I(_2929_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6965__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6957__A2 (.I(_2931_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A1 (.I(_2933_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6982__A2 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6964__A1 (.I(_2936_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6963__A2 (.I(_2937_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6969__A2 (.I(_2939_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6967__B2 (.I(_2941_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__A2 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6974__A1 (.I(_2947_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__B1 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__A2 (.I(_2948_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6997__A2 (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6976__B (.I(_2949_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6986__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6980__A2 (.I(_2953_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6990__B1 (.I(_2955_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6984__A2 (.I(_2957_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6988__B1 (.I(_2961_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7004__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7001__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6995__A2 (.I(_2967_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6998__A2 (.I(_2970_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7002__A2 (.I(_2973_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7016__A3 (.I(_2984_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A3 (.I(_2986_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7047__B (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7029__I (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7020__I (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7017__I (.I(_2988_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7026__I (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7025__I (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7021__I (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7019__I (.I(_2990_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A2 (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7043__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7032__I (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__B (.I(_2992_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7024__B (.I(_2995_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7031__A2 (.I(_2999_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7036__A2 (.I(_3004_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7040__A2 (.I(_3007_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7044__B (.I(_3011_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7048__B (.I(_3014_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7052__A2 (.I(_3016_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7056__A2 (.I(_3019_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7069__I (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7058__I (.I(_3021_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7068__A2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7066__A2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A2 (.I(_3022_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7070__I (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7060__I (.I(_3023_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7067__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7065__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7063__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7061__A2 (.I(_3024_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7077__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7075__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7073__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7071__A2 (.I(_3030_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7099__B2 (.I(_3040_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7088__A4 (.I(_3041_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7129__A3 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A1 (.I(_3046_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7095__A3 (.I(_3047_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7096__A2 (.I(_3049_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7123__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7098__A1 (.I(_3050_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A1 (.I(_3056_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7124__A2 (.I(_3057_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7110__A2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7109__B2 (.I(_3061_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7113__B2 (.I(_3064_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7121__A1 (.I(_3069_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A2 (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7134__C (.I(_3081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7156__A3 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7150__A3 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7144__A3 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7133__A2 (.I(_3084_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7154__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7148__A1 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7142__A2 (.I(_3092_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7171__A2 (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7165__I (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7160__I (.I(_3107_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7187__A2 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7184__B (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__B2 (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7161__B (.I(_3108_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7164__A2 (.I(_3109_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7181__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7180__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7175__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7166__A2 (.I(_3112_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7186__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7179__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7172__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7168__A1 (.I(_3114_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__S0 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3795__I (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__S1 (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3596__I (.I(_3131_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4136__I (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A1 (.I(_3133_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4746__I (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4139__C (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__A1 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3600__A2 (.I(_3135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4924__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4289__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A1 (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3602__I (.I(_3137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5192__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3753__A1 (.I(_3138_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A3 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A2 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3741__A1 (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3604__I (.I(_3139_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7015__A1 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A2 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4466__I (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3699__A1 (.I(_3140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6973__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5838__A2 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5836__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A1 (.I(_3141_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5443__I (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3689__A2 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3607__A2 (.I(_3142_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5206__I (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A2 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A1 (.I(_3147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5554__A1 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3614__A2 (.I(_3149_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3639__I (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3615__I (.I(_3150_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A2 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A1 (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3616__I (.I(_3151_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5136__I (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5057__B (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3700__I (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A1 (.I(_3152_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3743__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A2 (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3666__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3618__I (.I(_3153_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3633__I (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3631__A1 (.I(_3154_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5924__A2 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3721__A1 (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3670__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3620__I (.I(_3155_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5227__I (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A1 (.I(_3157_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3718__I (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A1 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A2 (.I(_3158_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4948__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A1 (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3624__I (.I(_3159_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3859__I (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3674__A2 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A1 (.I(_3160_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3869__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3637__I (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3628__A1 (.I(_3161_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3883__A2 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A3 (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3672__I (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3627__I (.I(_3162_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4110__I (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4067__B (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3982__A2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3629__A2 (.I(_3164_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A1 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4112__I (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A1 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3630__A3 (.I(_3165_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4791__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A2 (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3632__I (.I(_3167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7128__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5052__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3808__A1 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__A2 (.I(_3168_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5369__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4764__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A1 (.I(_3169_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4013__A1 (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3642__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3635__I (.I(_3170_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4492__A2 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A1 (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3636__I (.I(_3171_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5468__A1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5048__I (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A1 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A2 (.I(_3172_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A2 (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3638__I (.I(_3173_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5133__A3 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4993__A1 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A3 (.I(_3174_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4765__A1 (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3780__I (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3640__I (.I(_3175_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4777__A1 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4774__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4771__I (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3641__A4 (.I(_3176_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5010__I (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5007__A2 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A1 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A1 (.I(_3179_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4474__I (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3824__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3739__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A1 (.I(_3180_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5388__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4473__I (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3646__A2 (.I(_3181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6471__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5734__A1 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A2 (.I(_3184_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5654__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3954__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3763__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A1 (.I(_3185_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5650__A1 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4120__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3762__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3651__A2 (.I(_3186_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6644__I (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A2 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3652__A3 (.I(_3187_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4750__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A1 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3653__A2 (.I(_3188_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4800__A1 (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3654__B (.I(_3189_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__S (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3813__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3787__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3656__I (.I(_3191_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4296__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4293__A1 (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3785__S (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3658__I (.I(_3193_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__S (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__S (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3800__A1 (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3659__I (.I(_3194_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4743__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3717__I (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A1 (.I(_3195_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__S0 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A2 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__S0 (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3661__I (.I(_3196_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4489__I (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A2 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__S (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A1 (.I(_3197_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3922__A1 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3790__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3663__A2 (.I(_3198_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A2 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A2 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A2 (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3664__I (.I(_3199_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4752__A1 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3726__I (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3669__A2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3665__A2 (.I(_3200_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5038__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4483__A1 (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3667__I (.I(_3202_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5536__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4929__A2 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4801__A1 (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3668__I (.I(_3203_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5392__I (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5054__A1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A1 (.I(_3204_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4982__A1 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4488__I (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A1 (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3671__I (.I(_3206_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5612__I (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5474__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A1 (.I(_3207_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A1 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3860__A2 (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3673__I (.I(_3208_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5580__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4960__I (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4950__A1 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A2 (.I(_3209_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A3 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4930__A2 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4758__A2 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3676__A3 (.I(_3211_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6533__C (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5116__I (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5043__A2 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A3 (.I(_3212_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A3 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A3 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A3 (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3678__I (.I(_3213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5571__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A4 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A1 (.I(_3214_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4469__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A1 (.I(_3215_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A2 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4497__A2 (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4468__I (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3681__I (.I(_3216_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5444__A3 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4965__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3730__I (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3683__A1 (.I(_3218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__A2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5777__A2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4940__A2 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3684__A3 (.I(_3219_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5793__A1 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4763__A2 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3685__A2 (.I(_3220_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6701__A1 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6226__C (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6092__C (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3687__A4 (.I(_3222_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4754__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3846__A1 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3778__I (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3697__A2 (.I(_3227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6135__B2 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5649__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5504__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A1 (.I(_3228_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6184__B2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5652__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5506__A1 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3694__A2 (.I(_3229_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6685__A2 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6647__A2 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A3 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3695__A2 (.I(_3230_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6658__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5087__A2 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4983__I (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A1 (.I(_3236_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5842__B (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5708__B (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3703__A1 (.I(_3237_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3898__I (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A3 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3704__A1 (.I(_3239_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A1 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A2 (.I(_3241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A3 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3707__A2 (.I(_3242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7013__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5595__I (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4158__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3715__A1 (.I(_3244_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A2 (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3710__I (.I(_3245_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4256__A2 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4189__A1 (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__S (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3711__I (.I(_3246_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4180__I (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3713__A2 (.I(_3248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5795__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4775__A2 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3776__A1 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3716__A3 (.I(_3251_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5171__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4748__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3896__I (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A1 (.I(_3253_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5037__A1 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4964__A2 (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4740__I (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3719__I (.I(_3254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5481__B (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4797__A1 (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3767__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3720__I (.I(_3255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6464__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5090__I (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4480__A1 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A2 (.I(_3256_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4061__I (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3963__A2 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A1 (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3722__I (.I(_3257_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4329__A1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4323__A1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4257__A1 (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3724__I (.I(_3259_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4389__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4102__A2 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A1 (.I(_3261_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A3 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5042__A2 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5026__A3 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A3 (.I(_3262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3868__I (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3728__A1 (.I(_3263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5070__I (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A2 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3729__A4 (.I(_3264_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5385__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5356__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4968__I (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A1 (.I(_3266_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5814__A2 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5799__B (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4475__A1 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3733__A1 (.I(_3268_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5778__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5619__A3 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5607__A2 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3734__A3 (.I(_3269_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5858__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5518__I (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5455__A1 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3736__A2 (.I(_3271_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4885__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4744__A2 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A4 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3737__A4 (.I(_3272_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3959__I (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3751__A3 (.I(_3273_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5557__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5210__I (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4499__A2 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A1 (.I(_3274_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5044__I (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3740__A2 (.I(_3275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4155__I (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A1 (.I(_3276_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4159__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3907__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A1 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3742__A2 (.I(_3277_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4992__A2 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4760__A1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4481__I (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A1 (.I(_3279_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4015__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A1 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3745__A2 (.I(_3280_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3939__A1 (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3746__I (.I(_3281_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4780__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4354__A1 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4280__A1 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3747__A2 (.I(_3282_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A1 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5107__I (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4975__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3748__A2 (.I(_3283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4794__A2 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A3 (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3749__I (.I(_3284_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6463__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5046__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4773__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3750__A2 (.I(_3285_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__A1 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__A2 (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3752__I (.I(_3287_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4167__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4077__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A1 (.I(_3290_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5883__A2 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__I3 (.I(_3293_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4018__C (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3865__A2 (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3831__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3760__I (.I(_3295_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A1 (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3761__I (.I(_3296_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4014__I (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3854__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3765__A1 (.I(_3297_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A2 (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3766__I (.I(_3301_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6645__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6447__A2 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4789__A1 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3858__A1 (.I(_3302_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6472__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5579__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3897__I (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A1 (.I(_3303_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5751__A2 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5207__A2 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4470__A1 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3769__A2 (.I(_3304_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5733__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5556__A1 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A2 (.I(_3305_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6910__A1 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6723__B (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6681__I (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3772__A3 (.I(_3307_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4825__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3773__A1 (.I(_3308_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4309__A1 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4202__A1 (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3774__I (.I(_3309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7023__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6489__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5656__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__A1 (.I(_3311_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3949__I (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3843__I (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3777__I (.I(_3312_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6466__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5826__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5804__A1 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3779__A2 (.I(_3314_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4304__C (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__B (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__B (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3845__B (.I(_3315_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6474__A2 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5617__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5008__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3781__A1 (.I(_3316_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3944__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3915__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3841__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3782__I (.I(_3317_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7149__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7093__B (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6532__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A1 (.I(_3319_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6266__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3786__A2 (.I(_3321_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4208__S (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4133__I (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__S1 (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3788__I (.I(_3323_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__S (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4295__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4292__A1 (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3789__I (.I(_3324_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__S (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3799__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3793__A1 (.I(_3325_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4956__A1 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4433__A2 (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3794__B (.I(_3327_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4378__A3 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3801__A3 (.I(_3330_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__S0 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A2 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A1 (.I(_3331_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__C (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__C (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__C (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3797__A2 (.I(_3332_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4404__A1 (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3802__I (.I(_3337_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4411__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4403__A1 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4381__A2 (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3803__I (.I(_3338_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5159__A2 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4406__A1 (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3804__I (.I(_3339_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4888__A1 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A3 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4353__I (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__A2 (.I(_3340_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A1 (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3867__I (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3806__B (.I(_3341_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6457__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3844__A2 (.I(_3343_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4490__I (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4135__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4017__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3812__A1 (.I(_3346_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__S1 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__S (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__S1 (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3814__S (.I(_3349_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__I1 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3816__A2 (.I(_3350_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3910__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3818__I (.I(_3353_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A3 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A2 (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3819__I (.I(_3354_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4770__I (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3980__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3842__A2 (.I(_3355_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5247__A1 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5053__A2 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4954__A3 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A1 (.I(_3356_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5039__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4936__I (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3822__A2 (.I(_3357_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4762__I (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A2 (.I(_3358_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5513__A2 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4969__I (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A1 (.I(_3359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5798__A3 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3825__A2 (.I(_3360_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4467__A2 (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3826__I (.I(_3361_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5471__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5032__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5013__I (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3827__A3 (.I(_3362_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4859__A1 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3828__A2 (.I(_3363_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A1 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__A1 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A2 (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3832__I (.I(_3367_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A1 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3916__I (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3834__A2 (.I(_3369_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__A1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A3 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4768__A1 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3840__A2 (.I(_3370_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6679__A1 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A2 (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3837__I (.I(_3372_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5877__A2 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5179__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A1 (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3838__I (.I(_3373_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5884__A1 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5875__A1 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4757__I (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3839__A1 (.I(_3374_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6481__A3 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4782__A1 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3847__A2 (.I(_3382_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A1 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4033__I (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3912__B (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3853__A2 (.I(_3388_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6688__A2 (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3855__I (.I(_3390_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6649__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6445__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4785__A1 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3856__A2 (.I(_3391_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I0 (.I(_3394_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4078__I (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4068__I (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A1 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A1 (.I(_3395_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5025__A3 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4913__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4079__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3861__A2 (.I(_3396_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__B (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3966__A1 (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3892__I (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3862__I (.I(_3397_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4842__A1 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4400__A1 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4399__A1 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A1 (.I(_3398_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A1 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3877__A2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3866__A2 (.I(_3401_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4053__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3894__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A2 (.I(_3402_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__B (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3874__A1 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__A1 (.I(_3403_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4484__A2 (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__B (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3870__I (.I(_3405_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4103__I (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__A2 (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3879__A2 (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3871__A2 (.I(_3406_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4395__A1 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4183__C (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4092__A1 (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3873__B (.I(_3408_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7125__B (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__A1 (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A2 (.I(_3411_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5086__A1 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__A2 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3881__A2 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__A2 (.I(_3414_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4391__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4100__I (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A1 (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3880__B (.I(_3415_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4071__A1 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__B (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3886__A2 (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3884__I (.I(_3419_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4396__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4246__A2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4192__B2 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A1 (.I(_3420_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__B (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5077__A1 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A1 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3889__A2 (.I(_3421_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4933__A3 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3986__A1 (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3887__I (.I(_3422_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4398__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4397__C (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4337__A1 (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3888__B (.I(_3423_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4052__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3978__B (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3974__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3893__A2 (.I(_3427_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6450__A2 (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A1 (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4790__A1 (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__I1 (.I(_3431_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7143__A1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6548__A1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4799__A1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A1 (.I(_3432_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6462__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5861__A1 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5658__I (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A2 (.I(_3433_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5659__A2 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5469__A1 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5230__A4 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3899__A3 (.I(_3434_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3961__I (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3900__I (.I(_3435_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4234__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4164__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4074__A1 (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3901__S (.I(_3436_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7062__A1 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4438__A1 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3906__A2 (.I(_3437_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7059__B (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5531__I (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4435__B (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3903__B (.I(_3438_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4236__I (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3904__I (.I(_3439_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4166__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4076__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3992__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3905__A2 (.I(_3440_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4233__C (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4163__C (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3953__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3908__I (.I(_3442_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4057__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4049__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3956__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3913__A2 (.I(_3445_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6727__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6726__A2 (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3914__I (.I(_3448_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6496__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4818__A1 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3952__A2 (.I(_3449_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7104__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6503__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4813__A1 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3946__A2 (.I(_3451_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3920__A2 (.I(_3453_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4010__A1 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3923__A1 (.I(_3455_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4062__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3924__I (.I(_3458_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A2 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4122__A1 (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__B (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3925__I (.I(_3459_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7108__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4035__A2 (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3926__I (.I(_3460_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7033__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A3 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4812__A1 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3945__A2 (.I(_3461_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A1 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5998__A1 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A2 (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3928__I (.I(_3462_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5180__I (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5170__A2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__B2 (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3930__I (.I(_3464_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6689__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5941__A1 (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3931__I (.I(_3465_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5926__A1 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5125__I (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4811__A1 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3943__A1 (.I(_3466_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4196__A2 (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3936__I (.I(_3470_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4030__A2 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3972__A2 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3964__A2 (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3937__I (.I(_3471_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__B1 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A3 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3995__I (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3941__A1 (.I(_3472_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4409__A1 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4358__A1 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__A1 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3940__A2 (.I(_3473_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6499__A2 (.I(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5588__A4 (.I(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4810__A1 (.I(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3942__A2 (.I(_3476_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A2 (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4815__A1 (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4016__I0 (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3948__I (.I(_3482_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7028__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6493__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5670__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3950__A1 (.I(_3483_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3960__A2 (.I(_3487_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4425__A1 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4041__B (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__B (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3955__A2 (.I(_3489_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6720__A2 (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6719__A2 (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3957__I (.I(_3491_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6680__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6495__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4820__A1 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3958__A2 (.I(_3492_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3991__A1 (.I(_3495_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4235__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4165__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A1 (.I(_3496_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5672__I0 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3985__A1 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3981__A1 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3968__A1 (.I(_3502_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__C (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__B (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3987__A2 (.I(_3503_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5539__A1 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5244__A1 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4949__A3 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3970__A1 (.I(_3504_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4493__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4065__A1 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3977__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3971__A2 (.I(_3505_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5190__A2 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4392__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4255__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3976__A1 (.I(_3506_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A2 (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3975__A2 (.I(_3509_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3984__A1 (.I(_3511_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4184__I (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A1 (.I(_3512_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3979__A2 (.I(_3513_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3983__A2 (.I(_3514_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7106__A2 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3988__A2 (.I(_3522_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6498__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5073__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4821__A1 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3990__A2 (.I(_3524_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7064__A1 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4440__A1 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3993__A2 (.I(_3526_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5675__I (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A1 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4833__A1 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4027__A1 (.I(_3528_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7027__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6519__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5114__A1 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4026__A2 (.I(_3529_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3998__A2 (.I(_3530_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4082__A1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4001__A1 (.I(_3532_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4000__A2 (.I(_3533_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A2 (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4002__I (.I(_3535_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5587__A1 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A2 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4104__A2 (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4003__I (.I(_3536_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6549__A2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6535__B2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4230__A2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4025__A2 (.I(_3537_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6031__A2 (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4006__I (.I(_3539_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6753__A1 (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6752__B (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4007__I (.I(_3540_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__B (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B1 (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4008__I (.I(_3541_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A2 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A1 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4829__A1 (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4009__I (.I(_3542_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6748__A2 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6520__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5494__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4024__A1 (.I(_3543_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4028__I (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4011__I (.I(_3544_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4148__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4147__A4 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4034__A1 (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4012__I (.I(_3545_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5163__A2 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4847__A1 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4132__I (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4022__A1 (.I(_3546_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4934__A2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4357__B2 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A1 (.I(_3547_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7022__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6486__B2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5161__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4021__A2 (.I(_3548_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4221__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4020__A1 (.I(_3549_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4272__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4121__A2 (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4019__I (.I(_3552_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6522__A1 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5589__A1 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4830__A1 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4023__A2 (.I(_3556_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4069__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4046__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4045__A2 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4029__A3 (.I(_3562_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4118__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A1 (.I(_3563_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4039__A2 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4032__A2 (.I(_3564_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A2 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A1 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A1 (.I(_3566_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6760__A3 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6759__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4037__A2 (.I(_3570_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6729__A2 (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6514__A2 (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4835__A1 (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4038__A2 (.I(_3571_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4426__B2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4370__A1 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4200__B2 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4042__A1 (.I(_3574_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6722__A2 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6515__A2 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4836__A1 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4044__B1 (.I(_3577_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4075__A2 (.I(_3578_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4093__A2 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__A2 (.I(_3583_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5166__B2 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4417__A1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A1 (.I(_3584_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4054__B2 (.I(_3587_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4056__A2 (.I(_3589_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4094__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4089__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4058__A1 (.I(_3591_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4066__A2 (.I(_3593_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A1 (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6265__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5872__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5485__I (.I(\as2650.addr_buff[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6311__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5927__A1 (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5489__I (.I(\as2650.addr_buff[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6385__A3 (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5986__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5492__I (.I(\as2650.addr_buff[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6384__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6381__A1 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6055__B2 (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5496__I (.I(\as2650.addr_buff[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6996__B (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6421__A1 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6093__B2 (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5500__I (.I(\as2650.addr_buff[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3911__A1 (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3852__A1 (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3849__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3692__I (.I(\as2650.addr_buff[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4128__A2 (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3851__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3850__A2 (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3693__I (.I(\as2650.addr_buff[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6456__A1 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4051__A2 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3875__I (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A2 (.I(\as2650.carry ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5475__I (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5449__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3647__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3608__A1 (.I(\as2650.cycle[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4967__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3701__I (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A1 (.I(\as2650.halted ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5665__I0 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3891__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3864__A1 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3863__I0 (.I(\as2650.holding_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4107__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4081__I (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4080__A1 (.I(\as2650.holding_reg[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4334__I (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4330__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4316__A1 (.I(\as2650.holding_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7118__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4390__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4380__I (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4379__A1 (.I(\as2650.holding_reg[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3810__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__S0 (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3662__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3598__I (.I(\as2650.ins_reg[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3660__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3595__I (.I(\as2650.ins_reg[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3938__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A1 (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3634__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3622__I (.I(\as2650.ins_reg[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3727__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3623__I (.I(\as2650.ins_reg[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3882__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3744__A2 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3706__A1 (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3625__I (.I(\as2650.ins_reg[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7135__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6518__A1 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5165__B2 (.I(\as2650.overflow ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A3 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A1 (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4455__I (.I(\as2650.pc[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7006__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6417__A1 (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4572__I (.I(\as2650.pc[12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5975__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A1 (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5919__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4509__I (.I(\as2650.pc[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6051__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5969__A1 (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4514__I (.I(\as2650.pc[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A1 (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6025__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4520__I (.I(\as2650.pc[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A1 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6128__A2 (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6121__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4525__I (.I(\as2650.pc[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A1 (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4533__I (.I(\as2650.pc[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A1 (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4539__I (.I(\as2650.pc[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6257__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6211__A1 (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6207__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4544__I (.I(\as2650.pc[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A2 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6254__A1 (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4549__I (.I(\as2650.pc[8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6335__A1 (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6331__A1 (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6294__I (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4555__I (.I(\as2650.pc[9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7155__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5167__I (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5075__A1 (.I(\as2650.psl[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4050__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3876__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3805__A1 (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3783__I (.I(\as2650.psl[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3757__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3756__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3755__S (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3655__I (.I(\as2650.psl[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7100__B (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6561__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5169__A1 (.I(\as2650.psl[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7182__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6502__A1 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5181__B2 (.I(\as2650.psu[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7177__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6517__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__A1 (.I(\as2650.psu[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6530__I (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5187__B2 (.I(\as2650.psu[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5093__A3 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4783__A1 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3775__I (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3758__I0 (.I(\as2650.r0[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3947__I (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3815__A1 (.I(\as2650.r0[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3994__I (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3919__A1 (.I(\as2650.r0[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A4 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4848__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4154__I (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3997__A1 (.I(\as2650.r0[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A3 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4857__I (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4231__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4138__A1 (.I(\as2650.r0[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A2 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4984__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4278__I (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4210__A1 (.I(\as2650.r0[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5094__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4350__I (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4290__A1 (.I(\as2650.r0[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5155__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5095__B (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4421__I (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3784__A1 (.I(\as2650.r0[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6095__I0 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4237__A1 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4134__I1 (.I(\as2650.r123[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5289__I0 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3918__I1 (.I(\as2650.r123_2[1][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5291__I0 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3996__I1 (.I(\as2650.r123_2[1][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5938__I1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4822__I1 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3811__I3 (.I(\as2650.r123_2[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5997__I1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4840__I1 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3921__I3 (.I(\as2650.r123_2[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6044__I1 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4854__I1 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3999__I3 (.I(\as2650.r123_2[2][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6195__B2 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4720__A1 (.I(\as2650.stack[0][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__B2 (.I(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4726__I1 (.I(\as2650.stack[0][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__A1 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4696__A1 (.I(\as2650.stack[1][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__B2 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4676__A1 (.I(\as2650.stack[1][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__B2 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4679__A1 (.I(\as2650.stack[1][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__B2 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4682__A1 (.I(\as2650.stack[1][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6281__A1 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4686__I1 (.I(\as2650.stack[1][8] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6357__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4650__A1 (.I(\as2650.stack[2][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6395__C1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4652__A1 (.I(\as2650.stack[2][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6432__A1 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4654__A1 (.I(\as2650.stack[2][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5956__B2 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4628__A1 (.I(\as2650.stack[2][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6014__B2 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4630__A1 (.I(\as2650.stack[2][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6108__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4636__A1 (.I(\as2650.stack[2][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6152__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4638__A1 (.I(\as2650.stack[2][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6321__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4648__A1 (.I(\as2650.stack[2][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6356__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4612__A1 (.I(\as2650.stack[3][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6396__A1 (.I(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4614__A1 (.I(\as2650.stack[3][11] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6431__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4616__A1 (.I(\as2650.stack[3][12] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6106__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4598__A1 (.I(\as2650.stack[3][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6151__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4600__A1 (.I(\as2650.stack[3][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6194__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4602__A1 (.I(\as2650.stack[3][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6242__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4604__A1 (.I(\as2650.stack[3][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6322__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4610__A1 (.I(\as2650.stack[3][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6353__B2 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4565__A1 (.I(\as2650.stack[4][10] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__B2 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4531__A1 (.I(\as2650.stack[4][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__B2 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4537__A1 (.I(\as2650.stack[4][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__B2 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4547__A1 (.I(\as2650.stack[4][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6319__B2 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4560__A1 (.I(\as2650.stack[4][9] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5909__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5323__A1 (.I(\as2650.stack[5][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5325__A1 (.I(\as2650.stack[5][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6061__B2 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5329__A1 (.I(\as2650.stack[5][3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6103__B2 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5333__A1 (.I(\as2650.stack[5][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6147__B2 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5335__A1 (.I(\as2650.stack[5][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6191__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5337__A1 (.I(\as2650.stack[5][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6238__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5339__A1 (.I(\as2650.stack[5][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__B2 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5252__A1 (.I(\as2650.stack[6][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5960__C1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5254__A1 (.I(\as2650.stack[6][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6104__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5262__A1 (.I(\as2650.stack[6][4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6148__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5264__A1 (.I(\as2650.stack[6][5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6190__B2 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5266__A1 (.I(\as2650.stack[6][6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6239__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5268__A1 (.I(\as2650.stack[6][7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6600__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5911__A1 (.I(\as2650.stack[7][0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6602__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5961__A1 (.I(\as2650.stack[7][1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6604__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6011__A1 (.I(\as2650.stack[7][2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4656__A2 (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4577__I (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A2 (.I(\as2650.stack_ptr[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5409__A1 (.I(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4618__I (.I(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4578__A1 (.I(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4461__A1 (.I(\as2650.stack_ptr[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5901__A1 (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5411__A1 (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4465__I (.I(\as2650.stack_ptr[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7430__CLK (.I(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7274__CLK (.I(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7386__CLK (.I(clknet_leaf_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(wb_rst_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6697__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5937__A1 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5928__A2 (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3836__I (.I(net1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5939__A1 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5929__A2 (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3927__I (.I(net2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6030__A2 (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4004__I (.I(net3));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6027__A2 (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5185__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4143__I (.I(net4));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6166__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6081__A2 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5157__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4224__I (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6119__A2 (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4283__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6164__A2 (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4360__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6232__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4898__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__4413__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5839__C (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5001__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3902__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3702__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3603__A2 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output11_I (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output12_I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output13_I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output14_I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output15_I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output21_I (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5530__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output22_I (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5634__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5631__A1 (.I(net22));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output23_I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5604__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5601__A1 (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__3594__I (.I(net23));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output24_I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6576__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5178__I (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout52_I (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A2 (.I(net26));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output27_I (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6750__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6745__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6715__A1 (.I(net27));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_fanout51_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output31_I (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output32_I (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6881__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6865__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6842__A1 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output35_I (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6955__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6945__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6930__A1 (.I(net35));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output36_I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6977__I (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6971__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6956__A1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output37_I (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6993__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6991__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6979__A1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output38_I (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7009__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6994__A1 (.I(net38));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output41_I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7041__I (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output42_I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7045__I (.I(net42));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output43_I (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7051__A1 (.I(net43));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output44_I (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7055__A1 (.I(net44));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output45_I (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__5538__A1 (.I(net45));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6711__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output26_I (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6714__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__6676__A1 (.I(net52));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7336__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7198__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7301__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7199__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7191__CLK (.I(clknet_leaf_1_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7271__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7270__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7332__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7197__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7428__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7189__CLK (.I(clknet_leaf_2_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7304__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7337__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7433__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7429__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7190__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7333__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7339__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7338__CLK (.I(clknet_leaf_3_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7439__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7361__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7440__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7277__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7202__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7195__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7203__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7388__CLK (.I(clknet_leaf_6_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7284__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7449__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7362__CLK (.I(clknet_leaf_7_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7366__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7342__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7341__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7427__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7340__CLK (.I(clknet_leaf_14_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7424__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7425__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7420__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7423__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7426__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7422__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7421__CLK (.I(clknet_leaf_15_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7370__CLK (.I(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7348__CLK (.I(clknet_leaf_19_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7352__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7351__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7349__CLK (.I(clknet_leaf_21_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7385__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7373__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7376__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7330__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7329__CLK (.I(clknet_leaf_25_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7411__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7408__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7410__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7407__CLK (.I(clknet_leaf_27_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7417__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7415__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7414__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7416__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7418__CLK (.I(clknet_leaf_29_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7241__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7240__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7227__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7243__CLK (.I(clknet_leaf_31_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7214__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7269__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7217__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7215__CLK (.I(clknet_leaf_32_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7384__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7378__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7406__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7216__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7379__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7382__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7383__CLK (.I(clknet_leaf_33_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7405__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7404__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7296__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7297__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7299__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7298__CLK (.I(clknet_leaf_34_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7325__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7328__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7327__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7403__CLK (.I(clknet_leaf_35_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7238__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7211__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7213__CLK (.I(clknet_leaf_36_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7254__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7255__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7268__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7266__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7267__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7326__CLK (.I(clknet_leaf_37_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7253__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7224__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7225__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7229__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7242__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7230__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7228__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7256__CLK (.I(clknet_leaf_38_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7237__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7239__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7212__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7226__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7210__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7209__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7222__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7223__CLK (.I(clknet_leaf_39_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7250__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7249__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7263__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7251__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7236__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7235__CLK (.I(clknet_leaf_40_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7322__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7323__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7261__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7264__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7262__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7320__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7321__CLK (.I(clknet_leaf_42_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7265__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7324__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7402__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7295__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7397__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7290__CLK (.I(clknet_leaf_44_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7245__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7244__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7205__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7206__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7246__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7207__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7208__CLK (.I(clknet_leaf_48_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7287__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7288__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7394__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7395__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7396__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7219__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7220__CLK (.I(clknet_leaf_49_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7260__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7289__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7259__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7258__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7257__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7316__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7317__CLK (.I(clknet_leaf_50_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7372__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7363__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7437__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7436__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7444__CLK (.I(clknet_leaf_52_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7279__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7278__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7447__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7283__CLK (.I(clknet_leaf_53_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7446__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7442__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7448__CLK (.I(clknet_leaf_54_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7196__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7281__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7441__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7445__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7282__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7438__CLK (.I(clknet_leaf_60_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7306__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7307__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7305__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7204__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7275__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7276__CLK (.I(clknet_leaf_62_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7302__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7272__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7273__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7303__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7335__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7334__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7192__CLK (.I(clknet_leaf_64_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7357__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7355__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7356__CLK (.I(clknet_leaf_65_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0_0_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7358__CLK (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_65_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_64_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_63_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_10_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_2_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_1_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_0_wb_clk_i_I (.I(clknet_3_0_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_62_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_61_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_60_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_9_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_8_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_7_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_6_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7387__CLK (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_4_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_3_wb_clk_i_I (.I(clknet_3_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_17_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_16_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_15_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_14_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_13_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_12_wb_clk_i_I (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7393__CLK (.I(clknet_3_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_1_0_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7350__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_19_wb_clk_i_I (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7371__CLK (.I(clknet_3_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7443__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7314__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_57_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_56_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_54_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_53_wb_clk_i_I (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7280__CLK (.I(clknet_3_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_0_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_52_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_51_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_50_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_49_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_48_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_43_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__7374__CLK (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_24_wb_clk_i_I (.I(clknet_3_5_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_47_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_46_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_33_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_30_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_29_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_28_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_4_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_25_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_0_wb_clk_i_I (.I(clknet_3_6_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_45_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_44_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_42_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_41_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_40_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_39_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_38_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_37_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_36_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_35_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_34_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_32_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_31_wb_clk_i_I (.I(clknet_3_7_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_21_wb_clk_i_I (.I(clknet_opt_1_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_2_1_wb_clk_i_I (.I(clknet_opt_2_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_opt_3_1_wb_clk_i_I (.I(clknet_opt_3_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_leaf_27_wb_clk_i_I (.I(clknet_opt_4_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_1_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_1_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_1_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_1_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_1_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_1_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_1_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_2_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_2_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_2_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_2_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_2_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_2_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_2_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_3_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_3_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_3_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_3_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_3_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_3_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_3_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_4_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_4_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_4_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_4_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_4_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_4_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_4_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_5_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_5_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_5_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_5_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_6_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_6_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_6_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_6_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_6_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_7_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_7_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_7_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_7_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_8_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_8_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_8_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_8_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_8_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_9_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_9_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_9_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_9_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_10_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_10_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_10_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_10_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_10_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_11_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_11_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_11_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_11_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_12_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_12_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_12_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_12_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_12_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_13_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_13_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_13_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_13_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_14_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_14_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_14_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_14_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_14_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_15_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_15_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_15_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_15_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_16_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_16_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_16_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_16_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_16_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_17_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_17_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_17_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_17_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_18_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_18_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_18_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_18_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_18_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_19_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_19_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_19_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_19_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_20_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_20_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_20_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_20_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_20_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_21_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_21_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_21_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_21_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_22_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_22_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_22_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_22_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_22_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_23_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_23_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_23_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_23_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_23_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_23_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_23_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_24_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_24_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_24_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_24_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_24_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_24_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_25_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_25_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_25_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_25_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_25_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_25_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_25_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_26_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_26_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_26_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_26_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_26_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_27_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_27_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_27_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_27_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_28_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_28_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_28_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_28_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_28_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_29_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_29_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_29_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_29_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_30_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_30_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_30_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_30_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_30_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_31_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_31_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_31_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_31_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_32_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_32_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_32_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_32_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_32_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_33_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_33_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_33_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_33_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_34_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_34_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_34_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_34_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_34_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_35_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_35_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_35_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_35_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_36_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_36_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_36_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_36_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_36_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_37_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_37_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_37_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_37_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_38_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_38_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_38_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_38_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_38_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_39_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_39_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_39_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_39_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_40_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_40_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_40_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_40_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_40_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_41_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_41_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_41_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_41_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_42_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_42_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_42_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_42_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_42_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_42_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_42_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_43_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_43_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_43_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_43_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_43_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_43_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_43_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_44_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_44_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_44_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_44_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_44_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_44_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_44_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_45_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_45_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_45_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_45_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_45_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_45_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_45_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_46_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_46_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_46_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_46_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_46_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_46_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_46_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_47_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_47_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_47_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_47_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_47_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_47_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_47_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_48_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_48_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_48_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_48_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_48_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_48_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_48_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_49_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_49_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_49_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_49_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_49_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_49_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_49_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_50_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_50_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_50_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_50_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_50_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_50_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_50_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_51_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_51_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_51_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_51_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_51_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_51_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_52_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_52_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_52_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_52_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_52_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_52_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_52_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_53_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_53_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_53_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_53_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_53_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_53_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_53_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_54_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_54_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_54_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_54_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_54_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_54_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_54_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_55_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_55_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_55_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_55_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_55_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_55_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_56_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_56_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_56_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_56_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_56_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_56_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_56_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_57_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_57_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_57_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_57_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_57_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_57_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_57_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_58_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_58_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_58_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_58_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_58_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_58_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_58_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_59_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_59_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_59_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_59_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_59_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_59_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_59_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_60_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_60_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_60_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_60_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_60_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_60_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_60_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_61_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_61_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_61_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_61_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_61_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_61_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_61_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_62_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_62_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_62_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_62_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_62_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_62_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_62_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_27 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_63_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_63_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_63_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_63_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_63_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_63_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_63_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_64_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_64_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_64_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_64_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_64_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_64_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_64_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_65_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_65_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_65_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_65_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_65_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_65_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_65_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_66_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_66_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_66_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_66_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_66_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_66_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_66_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_67_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_67_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_67_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_67_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_67_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_67_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_67_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_68_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_68_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_68_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_68_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_68_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_68_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_68_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_69_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_69_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_69_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_69_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_69_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_69_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_69_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_70_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_70_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_70_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_70_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_70_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_70_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_70_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_71_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_71_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_71_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_71_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_71_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_71_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_71_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_72_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_72_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_72_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_72_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_72_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_72_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_72_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_73_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_73_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_73_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_73_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_73_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_73_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_74_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_74_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_74_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_74_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_74_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_74_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_74_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_75_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_75_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_75_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_75_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_75_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_75_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_76_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_76_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_76_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_76_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_76_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_76_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_76_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_77_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_77_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_77_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_77_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_77_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_77_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_78_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_78_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_78_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_78_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_78_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_78_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_78_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_79_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_79_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_79_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_79_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_79_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_79_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_79_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_80_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_80_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_80_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_80_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_80_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_80_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_80_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_81_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_81_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_81_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_81_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_81_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_81_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_81_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_82_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_82_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_82_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_82_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_82_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_82_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_82_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_83_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_83_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_83_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_83_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_83_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_83_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_83_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_84_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_84_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_84_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_84_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_84_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_84_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_84_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_85_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_85_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_85_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_85_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_85_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_85_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_85_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_355 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_86_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_86_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_86_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_86_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_86_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_86_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_86_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_21 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_87_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_87_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_87_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_87_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_87_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_87_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_87_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_88_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_88_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_88_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_88_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_88_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_88_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_88_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_89_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_89_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_89_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_89_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_89_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_89_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_90_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_90_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_90_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_90_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_90_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_90_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_90_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_91_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_91_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_91_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_91_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_91_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_91_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_23 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_25 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_474 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_92_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_92_1375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_92_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_92_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_92_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_92_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_92_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_93_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_93_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_93_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_93_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_93_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_93_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_93_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_574 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_94_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_94_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_94_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_94_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_94_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_94_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_94_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_31 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_95_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_95_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_95_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_95_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_95_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_95_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_95_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_96_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_96_1372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1380 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_96_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_96_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_96_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_96_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_96_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_604 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_97_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_97_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_97_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_97_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_97_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_97_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_97_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_514 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_98_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_98_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_98_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_98_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_98_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_98_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_98_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_390 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_615 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_99_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_99_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1035 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_99_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_99_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_99_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_99_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_99_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_100_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_100_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_100_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_100_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_100_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_100_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_100_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_101_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_101_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_101_1341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_101_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_101_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_101_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_101_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_19 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_102_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_102_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_102_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_102_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_102_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_102_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_102_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_103_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_103_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_103_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_103_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_103_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_103_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_103_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_104_1369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_104_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_104_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_104_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_104_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_104_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_104_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_17 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_596 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_105_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_105_1365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_105_1417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_105_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_105_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_105_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_105_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_7 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_11 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_15 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_106_1373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_106_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_106_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_106_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_106_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_106_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_106_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_107_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_626 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_107_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_107_1418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_107_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_107_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_107_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_107_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_108_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1065 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1083 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_108_1381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_108_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_108_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_108_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_108_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_108_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_109_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1116 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_109_1336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_109_1340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_109_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_109_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_109_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_109_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_429 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_711 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_110_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1001 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_110_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_110_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_110_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_110_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_110_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_110_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_111_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_111_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_111_1347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_111_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_111_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_111_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_111_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_451 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_836 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_980 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1090 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_112_1370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_112_1382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_112_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_112_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_112_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_112_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_112_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1086 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1088 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1268 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1284 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_113_1288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_113_1298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_113_1346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_113_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_113_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_113_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_113_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_427 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_114_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_822 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_923 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_114_1239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_114_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_114_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_114_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_114_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_114_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_20 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_115_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_661 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_115_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_115_1199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_115_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_115_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_115_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_115_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_498 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_575 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_879 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1071 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_116_1180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_116_1233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_116_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_116_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_116_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_116_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_116_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_464 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1007 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_117_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_117_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_117_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_117_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_117_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_117_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_117_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_442 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_453 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_701 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_997 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_118_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_118_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_118_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_118_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_118_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_118_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_118_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_538 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_544 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_616 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1091 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_119_1159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_119_1163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_119_1195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_119_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_119_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_119_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_119_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_280 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_284 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_549 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_120_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1045 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1073 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_120_1147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_120_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_120_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_120_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_120_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_120_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_414 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_468 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_540 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_121_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1029 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1037 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1039 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_121_1151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_121_1155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_121_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_121_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_121_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_121_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_537 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_651 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_671 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_828 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_122_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_984 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1008 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1068 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1096 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_122_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_122_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_122_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_122_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_122_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_122_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_123_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_965 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1002 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1006 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_123_1018 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1082 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_123_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_123_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_123_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_123_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_123_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_441 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_581 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_645 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_852 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1000 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1010 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1048 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1056 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_124_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1089 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_124_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_124_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_124_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_124_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_124_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_124_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_323 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_125_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_434 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_478 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_558 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_832 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_888 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_125_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_939 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_125_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_125_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_125_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_125_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_125_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_431 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_438 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_708 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_714 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_126_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1059 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1072 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1076 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1098 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_126_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_126_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_126_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_126_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_126_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_126_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_465 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_536 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_560 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_633 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_773 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_848 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_862 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_964 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_972 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1053 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1061 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1085 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_127_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_127_1193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_127_1205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_127_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_127_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_127_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_127_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_477 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_497 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_500 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_508 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_858 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_946 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1004 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1016 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1046 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_128_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_128_1123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_128_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_128_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_128_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_128_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_128_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_361 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_394 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_505 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_509 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_622 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_678 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_696 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_764 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_129_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1047 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1092 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_129_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_129_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_129_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_129_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_129_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_426 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_548 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_685 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_771 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_785 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_806 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_860 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_924 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_986 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1041 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1055 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1066 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1080 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1140 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_130_1160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_130_1168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_130_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_130_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_130_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_130_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_130_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_281 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_423 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_512 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_516 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_532 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_590 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_618 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_674 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_131_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_720 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_748 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_899 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_953 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_961 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_985 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1036 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1040 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1043 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_131_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1062 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_131_1133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_131_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_131_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_131_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_131_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_367 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_501 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_504 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_520 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_556 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_569 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_594 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_639 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_650 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_787 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_825 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_864 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_868 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_872 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_876 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_916 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_962 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_988 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1012 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1024 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1044 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1058 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1074 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1078 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1121 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1125 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_132_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_132_1169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_132_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_132_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_132_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_132_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_132_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_182 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_133_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_350 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_398 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_415 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_519 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_591 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_680 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_684 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_728 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_732 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_746 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_846 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_849 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_857 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_914 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_952 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_956 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_966 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_970 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_974 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_978 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1030 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1038 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1042 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1051 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1057 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1075 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1079 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1094 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_133_1107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_133_1127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_133_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_133_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_133_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_133_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_395 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_435 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_445 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_449 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_483 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_529 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_568 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_595 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_612 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_662 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_679 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_692 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_697 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_700 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_704 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_736 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_740 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_793 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_795 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_841 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_870 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_880 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_884 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_898 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_902 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_928 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_950 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_977 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_134_981 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1034 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1050 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1054 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1093 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_134_1097 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_134_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_134_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_134_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_134_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_134_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_430 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_446 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_480 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_513 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_517 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_521 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_561 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_592 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_599 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_630 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_637 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_653 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_655 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_658 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_670 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_688 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_693 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_731 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_753 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_761 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_802 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_805 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_819 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_829 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_833 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_856 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_866 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_890 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_894 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_135_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_931 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_949 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_959 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_969 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_973 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_989 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1005 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1020 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_135_1032 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1070 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_135_1134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_135_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_135_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_135_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_135_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_409 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_443 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_450 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_541 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_545 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_553 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_578 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_586 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_613 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_617 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_727 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_751 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_768 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_774 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_781 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_812 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_136_834 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_900 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_911 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_915 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_930 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_936 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_940 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_995 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_136_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1025 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_136_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_136_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_136_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_136_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_136_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_421 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_455 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_467 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_473 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_506 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_522 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_539 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_579 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_583 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_587 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_603 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_619 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_627 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_647 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_663 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_681 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_683 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_705 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_739 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_767 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_790 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_810 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_816 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_820 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_824 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_844 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_847 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_875 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_883 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_887 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_891 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_895 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_910 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_918 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_922 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_934 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_948 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_137_983 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_137_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_137_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_137_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_137_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_137_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_258 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_371 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_385 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_432 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_436 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_459 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_470 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_502 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_518 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_526 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_530 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_566 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_582 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_588 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_598 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_621 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_625 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_628 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_640 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_648 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_652 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_665 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_690 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_694 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_713 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_725 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_754 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_758 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_770 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_778 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_789 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_797 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_801 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_809 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_813 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_823 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_855 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_903 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_907 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_938 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_942 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_994 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_998 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_138_1014 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1022 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_138_1026 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1028 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_138_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_138_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_138_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_138_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_138_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_292 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_376 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_388 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_396 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_454 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_471 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_475 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_495 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_503 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_511 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_525 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_535 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_543 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_577 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_585 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_610 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_614 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_620 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_624 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_636 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_666 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_669 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_677 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_687 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_695 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_735 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_743 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_750 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_760 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_762 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_775 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_786 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_791 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_826 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_139_830 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_838 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_840 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_932 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_944 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_954 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_958 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_990 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_999 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_139_1063 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_139_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_139_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_139_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_139_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_370 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_386 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_401 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_412 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_487 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_491 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_546 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_584 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_600 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_611 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_623 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_631 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_642 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_646 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_654 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_656 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_659 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_689 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_703 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_719 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_723 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_730 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_752 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_756 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_766 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_776 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_788 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_794 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_798 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_814 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_827 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_835 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_853 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_861 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_865 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_878 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_882 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_886 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_908 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_917 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_945 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1011 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_140_1015 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1023 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_140_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_140_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_140_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_140_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_140_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_140_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_283 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_407 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_444 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_452 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_462 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_466 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_488 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_510 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_542 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_552 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_555 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_565 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_141_573 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_634 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_657 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_698 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_716 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_729 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_745 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_792 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_800 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_831 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_843 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_845 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_851 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_881 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_141_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_893 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_906 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_913 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_919 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_968 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_976 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_141_992 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_141_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_141_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_141_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_141_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_191 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_389 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_424 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_440 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_448 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_456 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_460 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_463 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_479 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_482 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_524 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_534 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_550 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_554 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_571 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_605 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_609 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_664 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_673 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_676 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_706 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_710 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_718 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_722 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_726 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_734 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_744 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_747 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_755 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_759 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_763 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_815 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_821 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_837 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_885 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_889 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_897 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_904 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_920 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_926 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_957 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_960 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_963 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_971 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1003 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_142_1019 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_142_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1031 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1095 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1099 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1315 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1386 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1450 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1454 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_142_1457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1521 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1525 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_142_1528 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_142_1560 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_142_1576 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_142_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_5 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_141 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_340 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_360 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_392 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_420 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_428 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_458 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_490 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_494 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_496 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_499 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_533 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_570 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_602 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_606 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_608 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_638 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_641 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_644 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_660 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_668 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_672 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_675 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_707 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_709 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_712 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_715 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_724 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_738 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_742 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_749 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_780 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_783 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_796 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_804 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_808 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_818 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_863 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_869 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_873 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_143_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_921 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_925 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_929 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_933 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_937 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_941 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_143_955 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_143_991 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_993 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_996 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1067 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1206 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1277 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1280 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1415 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1486 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1490 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_143_1493 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1557 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1561 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_143_1564 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_143_1572 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_143_1580 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_9 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_13 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_29 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_369 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_422 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_425 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_433 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_439 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_457 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_472 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_476 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_481 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_485 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_492 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_515 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_527 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_551 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_559 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_562 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_589 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_593 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_597 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_601 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_607 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_629 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_632 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_635 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_643 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_649 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_667 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_682 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_686 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_691 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_699 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_702 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_717 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_721 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_733 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_737 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_741 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_757 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_765 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_769 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_772 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_777 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_779 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_782 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_784 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_799 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_803 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_807 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_811 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_817 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_839 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_842 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_850 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_854 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_859 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_867 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_871 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_874 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_877 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_892 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_896 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_901 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_905 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_909 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_912 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_927 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_935 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_943 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_947 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_951 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_967 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_975 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_979 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_982 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_987 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1009 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1013 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1017 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1021 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1027 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1033 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1049 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1052 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1060 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1064 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1069 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1077 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1081 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1084 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1087 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1122 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1137 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1145 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1153 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1227 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1259 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1270 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1293 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1297 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1332 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1353 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1357 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1367 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1371 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1399 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1402 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1407 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1437 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1441 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1447 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1455 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1461 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1469 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1472 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1480 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1484 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1489 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1497 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1503 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1507 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1523 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_144_1531 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1539 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_144_1542 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_144_1547 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1563 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1567 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_144_1573 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_144_1577 ();
 assign io_oeb[10] = net54;
 assign io_oeb[11] = net55;
 assign io_oeb[12] = net56;
 assign io_oeb[13] = net57;
 assign io_oeb[14] = net58;
 assign io_oeb[15] = net59;
 assign io_oeb[16] = net60;
 assign io_oeb[17] = net61;
 assign io_oeb[18] = net62;
 assign io_oeb[19] = net63;
 assign io_oeb[20] = net64;
 assign io_oeb[21] = net65;
 assign io_oeb[22] = net66;
 assign io_oeb[23] = net67;
 assign io_oeb[24] = net68;
 assign io_oeb[25] = net69;
 assign io_oeb[26] = net70;
 assign io_oeb[27] = net71;
 assign io_oeb[28] = net72;
 assign io_oeb[29] = net73;
 assign io_oeb[30] = net74;
 assign io_oeb[31] = net75;
 assign io_oeb[32] = net76;
 assign io_oeb[33] = net77;
 assign io_oeb[34] = net78;
 assign io_oeb[35] = net79;
 assign io_oeb[36] = net80;
 assign io_oeb[37] = net81;
 assign io_oeb[8] = net93;
 assign io_oeb[9] = net53;
 assign io_out[28] = net83;
 assign io_out[29] = net84;
 assign io_out[30] = net85;
 assign io_out[31] = net86;
 assign io_out[32] = net87;
 assign io_out[33] = net88;
 assign io_out[34] = net89;
 assign io_out[35] = net90;
 assign io_out[36] = net91;
 assign io_out[37] = net92;
 assign io_out[8] = net82;
endmodule

