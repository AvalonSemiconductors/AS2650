VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO wrapped_as2650
  CLASS BLOCK ;
  FOREIGN wrapped_as2650 ;
  ORIGIN 0.000 0.000 ;
  SIZE 1050.000 BY 700.000 ;
  PIN RAM_end_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 409.920 4.000 410.480 ;
    END
  END RAM_end_addr[0]
  PIN RAM_end_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 477.120 4.000 477.680 ;
    END
  END RAM_end_addr[10]
  PIN RAM_end_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 483.840 4.000 484.400 ;
    END
  END RAM_end_addr[11]
  PIN RAM_end_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 490.560 4.000 491.120 ;
    END
  END RAM_end_addr[12]
  PIN RAM_end_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 497.280 4.000 497.840 ;
    END
  END RAM_end_addr[13]
  PIN RAM_end_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 504.000 4.000 504.560 ;
    END
  END RAM_end_addr[14]
  PIN RAM_end_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 510.720 4.000 511.280 ;
    END
  END RAM_end_addr[15]
  PIN RAM_end_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 416.640 4.000 417.200 ;
    END
  END RAM_end_addr[1]
  PIN RAM_end_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 423.360 4.000 423.920 ;
    END
  END RAM_end_addr[2]
  PIN RAM_end_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 430.080 4.000 430.640 ;
    END
  END RAM_end_addr[3]
  PIN RAM_end_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 436.800 4.000 437.360 ;
    END
  END RAM_end_addr[4]
  PIN RAM_end_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 443.520 4.000 444.080 ;
    END
  END RAM_end_addr[5]
  PIN RAM_end_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 450.240 4.000 450.800 ;
    END
  END RAM_end_addr[6]
  PIN RAM_end_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 456.960 4.000 457.520 ;
    END
  END RAM_end_addr[7]
  PIN RAM_end_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 463.680 4.000 464.240 ;
    END
  END RAM_end_addr[8]
  PIN RAM_end_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 470.400 4.000 470.960 ;
    END
  END RAM_end_addr[9]
  PIN RAM_start_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 275.520 4.000 276.080 ;
    END
  END RAM_start_addr[0]
  PIN RAM_start_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.720 4.000 343.280 ;
    END
  END RAM_start_addr[10]
  PIN RAM_start_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 349.440 4.000 350.000 ;
    END
  END RAM_start_addr[11]
  PIN RAM_start_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 356.160 4.000 356.720 ;
    END
  END RAM_start_addr[12]
  PIN RAM_start_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.880 4.000 363.440 ;
    END
  END RAM_start_addr[13]
  PIN RAM_start_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 369.600 4.000 370.160 ;
    END
  END RAM_start_addr[14]
  PIN RAM_start_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 376.320 4.000 376.880 ;
    END
  END RAM_start_addr[15]
  PIN RAM_start_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 282.240 4.000 282.800 ;
    END
  END RAM_start_addr[1]
  PIN RAM_start_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.960 4.000 289.520 ;
    END
  END RAM_start_addr[2]
  PIN RAM_start_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.680 4.000 296.240 ;
    END
  END RAM_start_addr[3]
  PIN RAM_start_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.400 4.000 302.960 ;
    END
  END RAM_start_addr[4]
  PIN RAM_start_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 309.120 4.000 309.680 ;
    END
  END RAM_start_addr[5]
  PIN RAM_start_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.840 4.000 316.400 ;
    END
  END RAM_start_addr[6]
  PIN RAM_start_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 322.560 4.000 323.120 ;
    END
  END RAM_start_addr[7]
  PIN RAM_start_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 329.280 4.000 329.840 ;
    END
  END RAM_start_addr[8]
  PIN RAM_start_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 336.000 4.000 336.560 ;
    END
  END RAM_start_addr[9]
  PIN WEb_ram
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 665.280 696.000 665.840 700.000 ;
    END
  END WEb_ram
  PIN boot_rom_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 403.200 4.000 403.760 ;
    END
  END boot_rom_en
  PIN bus_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 477.120 696.000 477.680 700.000 ;
    END
  END bus_addr[0]
  PIN bus_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 490.560 696.000 491.120 700.000 ;
    END
  END bus_addr[1]
  PIN bus_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 504.000 696.000 504.560 700.000 ;
    END
  END bus_addr[2]
  PIN bus_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 517.440 696.000 518.000 700.000 ;
    END
  END bus_addr[3]
  PIN bus_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 530.880 696.000 531.440 700.000 ;
    END
  END bus_addr[4]
  PIN bus_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 544.320 696.000 544.880 700.000 ;
    END
  END bus_addr[5]
  PIN bus_cyc
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 463.680 696.000 464.240 700.000 ;
    END
  END bus_cyc
  PIN bus_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 356.160 696.000 356.720 700.000 ;
    END
  END bus_data_out[0]
  PIN bus_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 369.600 696.000 370.160 700.000 ;
    END
  END bus_data_out[1]
  PIN bus_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 383.040 696.000 383.600 700.000 ;
    END
  END bus_data_out[2]
  PIN bus_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 396.480 696.000 397.040 700.000 ;
    END
  END bus_data_out[3]
  PIN bus_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 409.920 696.000 410.480 700.000 ;
    END
  END bus_data_out[4]
  PIN bus_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 423.360 696.000 423.920 700.000 ;
    END
  END bus_data_out[5]
  PIN bus_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 436.800 696.000 437.360 700.000 ;
    END
  END bus_data_out[6]
  PIN bus_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 450.240 696.000 450.800 700.000 ;
    END
  END bus_data_out[7]
  PIN bus_in_gpios[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 440.160 1050.000 440.720 ;
    END
  END bus_in_gpios[0]
  PIN bus_in_gpios[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 446.880 1050.000 447.440 ;
    END
  END bus_in_gpios[1]
  PIN bus_in_gpios[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 453.600 1050.000 454.160 ;
    END
  END bus_in_gpios[2]
  PIN bus_in_gpios[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 460.320 1050.000 460.880 ;
    END
  END bus_in_gpios[3]
  PIN bus_in_gpios[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 467.040 1050.000 467.600 ;
    END
  END bus_in_gpios[4]
  PIN bus_in_gpios[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 473.760 1050.000 474.320 ;
    END
  END bus_in_gpios[5]
  PIN bus_in_gpios[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 480.480 1050.000 481.040 ;
    END
  END bus_in_gpios[6]
  PIN bus_in_gpios[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 487.200 1050.000 487.760 ;
    END
  END bus_in_gpios[7]
  PIN bus_in_serial_ports[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 557.760 696.000 558.320 700.000 ;
    END
  END bus_in_serial_ports[0]
  PIN bus_in_serial_ports[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 571.200 696.000 571.760 700.000 ;
    END
  END bus_in_serial_ports[1]
  PIN bus_in_serial_ports[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 584.640 696.000 585.200 700.000 ;
    END
  END bus_in_serial_ports[2]
  PIN bus_in_serial_ports[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 598.080 696.000 598.640 700.000 ;
    END
  END bus_in_serial_ports[3]
  PIN bus_in_serial_ports[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 611.520 696.000 612.080 700.000 ;
    END
  END bus_in_serial_ports[4]
  PIN bus_in_serial_ports[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 624.960 696.000 625.520 700.000 ;
    END
  END bus_in_serial_ports[5]
  PIN bus_in_serial_ports[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 638.400 696.000 638.960 700.000 ;
    END
  END bus_in_serial_ports[6]
  PIN bus_in_serial_ports[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 651.840 696.000 652.400 700.000 ;
    END
  END bus_in_serial_ports[7]
  PIN bus_in_sid[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 507.360 1050.000 507.920 ;
    END
  END bus_in_sid[0]
  PIN bus_in_sid[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 514.080 1050.000 514.640 ;
    END
  END bus_in_sid[1]
  PIN bus_in_sid[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 520.800 1050.000 521.360 ;
    END
  END bus_in_sid[2]
  PIN bus_in_sid[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 527.520 1050.000 528.080 ;
    END
  END bus_in_sid[3]
  PIN bus_in_sid[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 534.240 1050.000 534.800 ;
    END
  END bus_in_sid[4]
  PIN bus_in_sid[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 540.960 1050.000 541.520 ;
    END
  END bus_in_sid[5]
  PIN bus_in_sid[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 547.680 1050.000 548.240 ;
    END
  END bus_in_sid[6]
  PIN bus_in_sid[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 554.400 1050.000 554.960 ;
    END
  END bus_in_sid[7]
  PIN bus_in_timers[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 947.520 696.000 948.080 700.000 ;
    END
  END bus_in_timers[0]
  PIN bus_in_timers[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 960.960 696.000 961.520 700.000 ;
    END
  END bus_in_timers[1]
  PIN bus_in_timers[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 974.400 696.000 974.960 700.000 ;
    END
  END bus_in_timers[2]
  PIN bus_in_timers[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 987.840 696.000 988.400 700.000 ;
    END
  END bus_in_timers[3]
  PIN bus_in_timers[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1001.280 696.000 1001.840 700.000 ;
    END
  END bus_in_timers[4]
  PIN bus_in_timers[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1014.720 696.000 1015.280 700.000 ;
    END
  END bus_in_timers[5]
  PIN bus_in_timers[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1028.160 696.000 1028.720 700.000 ;
    END
  END bus_in_timers[6]
  PIN bus_in_timers[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1041.600 696.000 1042.160 700.000 ;
    END
  END bus_in_timers[7]
  PIN bus_we_gpios
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 433.440 1050.000 434.000 ;
    END
  END bus_we_gpios
  PIN bus_we_serial_ports
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 934.080 696.000 934.640 700.000 ;
    END
  END bus_we_serial_ports
  PIN bus_we_sid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 500.640 1050.000 501.200 ;
    END
  END bus_we_sid
  PIN bus_we_timers
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 920.640 696.000 921.200 700.000 ;
    END
  END bus_we_timers
  PIN cs_port[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 383.040 4.000 383.600 ;
    END
  END cs_port[0]
  PIN cs_port[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.760 4.000 390.320 ;
    END
  END cs_port[1]
  PIN cs_port[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 396.480 4.000 397.040 ;
    END
  END cs_port[2]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.102000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 6.720 696.000 7.280 700.000 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 141.120 696.000 141.680 700.000 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 154.560 696.000 155.120 700.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 168.000 696.000 168.560 700.000 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 181.440 696.000 182.000 700.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 194.880 696.000 195.440 700.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 208.320 696.000 208.880 700.000 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 221.760 696.000 222.320 700.000 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 235.200 696.000 235.760 700.000 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 248.640 696.000 249.200 700.000 ;
    END
  END io_in[18]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 20.160 696.000 20.720 700.000 ;
    END
  END io_in[1]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 33.600 696.000 34.160 700.000 ;
    END
  END io_in[2]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 47.040 696.000 47.600 700.000 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.183000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 60.480 696.000 61.040 700.000 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.920 696.000 74.480 700.000 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 87.360 696.000 87.920 700.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 696.000 101.360 700.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 696.000 114.800 700.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 127.680 696.000 128.240 700.000 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.840 4.000 148.400 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 215.040 4.000 215.600 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.760 4.000 222.320 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 228.480 4.000 229.040 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 235.200 4.000 235.760 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.920 4.000 242.480 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.640 4.000 249.200 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 255.360 4.000 255.920 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.080 4.000 262.640 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.800 4.000 269.360 ;
    END
  END io_oeb[18]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 154.560 4.000 155.120 ;
    END
  END io_oeb[1]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 161.280 4.000 161.840 ;
    END
  END io_oeb[2]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 168.000 4.000 168.560 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.720 4.000 175.280 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 181.440 4.000 182.000 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 188.160 4.000 188.720 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.880 4.000 195.440 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 201.600 4.000 202.160 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 208.320 4.000 208.880 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 20.160 4.000 20.720 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 87.360 4.000 87.920 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.800 4.000 101.360 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 107.520 4.000 108.080 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.960 4.000 121.520 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.897600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.400 4.000 134.960 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 141.120 4.000 141.680 ;
    END
  END io_out[18]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 26.880 4.000 27.440 ;
    END
  END io_out[1]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 33.600 4.000 34.160 ;
    END
  END io_out[2]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 40.320 4.000 40.880 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 47.040 4.000 47.600 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.760 4.000 54.320 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 60.480 4.000 61.040 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 67.200 4.000 67.760 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.920 4.000 74.480 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.640 4.000 81.200 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 413.280 1050.000 413.840 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 420.000 1050.000 420.560 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 426.720 1050.000 427.280 ;
    END
  END irq[2]
  PIN irqs[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 262.080 696.000 262.640 700.000 ;
    END
  END irqs[0]
  PIN irqs[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 275.520 696.000 276.080 700.000 ;
    END
  END irqs[1]
  PIN irqs[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 288.960 696.000 289.520 700.000 ;
    END
  END irqs[2]
  PIN irqs[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 302.400 696.000 302.960 700.000 ;
    END
  END irqs[3]
  PIN irqs[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 315.840 696.000 316.400 700.000 ;
    END
  END irqs[4]
  PIN irqs[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 329.280 696.000 329.840 700.000 ;
    END
  END irqs[5]
  PIN irqs[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 342.720 696.000 343.280 700.000 ;
    END
  END irqs[6]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 36.960 1050.000 37.520 ;
    END
  END la_data_out[0]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 104.160 1050.000 104.720 ;
    END
  END la_data_out[10]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 110.880 1050.000 111.440 ;
    END
  END la_data_out[11]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 117.600 1050.000 118.160 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 124.320 1050.000 124.880 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 131.040 1050.000 131.600 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 137.760 1050.000 138.320 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 144.480 1050.000 145.040 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 151.200 1050.000 151.760 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 157.920 1050.000 158.480 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 164.640 1050.000 165.200 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 43.680 1050.000 44.240 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 171.360 1050.000 171.920 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 178.080 1050.000 178.640 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 184.800 1050.000 185.360 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 191.520 1050.000 192.080 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 198.240 1050.000 198.800 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 204.960 1050.000 205.520 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 211.680 1050.000 212.240 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 218.400 1050.000 218.960 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 225.120 1050.000 225.680 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 231.840 1050.000 232.400 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 50.400 1050.000 50.960 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 238.560 1050.000 239.120 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 245.280 1050.000 245.840 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 252.000 1050.000 252.560 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 258.720 1050.000 259.280 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 265.440 1050.000 266.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 272.160 1050.000 272.720 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 278.880 1050.000 279.440 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 285.600 1050.000 286.160 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 292.320 1050.000 292.880 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 299.040 1050.000 299.600 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 57.120 1050.000 57.680 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 305.760 1050.000 306.320 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 312.480 1050.000 313.040 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 319.200 1050.000 319.760 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 325.920 1050.000 326.480 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 332.640 1050.000 333.200 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 339.360 1050.000 339.920 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 346.080 1050.000 346.640 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 352.800 1050.000 353.360 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 359.520 1050.000 360.080 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 366.240 1050.000 366.800 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 63.840 1050.000 64.400 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 372.960 1050.000 373.520 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 379.680 1050.000 380.240 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 386.400 1050.000 386.960 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 393.120 1050.000 393.680 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 399.840 1050.000 400.400 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.536800 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 406.560 1050.000 407.120 ;
    END
  END la_data_out[55]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 70.560 1050.000 71.120 ;
    END
  END la_data_out[5]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 77.280 1050.000 77.840 ;
    END
  END la_data_out[6]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 84.000 1050.000 84.560 ;
    END
  END la_data_out[7]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 90.720 1050.000 91.280 ;
    END
  END la_data_out[8]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 97.440 1050.000 98.000 ;
    END
  END la_data_out[9]
  PIN last_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 705.600 696.000 706.160 700.000 ;
    END
  END last_addr[0]
  PIN last_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 840.000 696.000 840.560 700.000 ;
    END
  END last_addr[10]
  PIN last_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 853.440 696.000 854.000 700.000 ;
    END
  END last_addr[11]
  PIN last_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 866.880 696.000 867.440 700.000 ;
    END
  END last_addr[12]
  PIN last_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 880.320 696.000 880.880 700.000 ;
    END
  END last_addr[13]
  PIN last_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 893.760 696.000 894.320 700.000 ;
    END
  END last_addr[14]
  PIN last_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 907.200 696.000 907.760 700.000 ;
    END
  END last_addr[15]
  PIN last_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 719.040 696.000 719.600 700.000 ;
    END
  END last_addr[1]
  PIN last_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 732.480 696.000 733.040 700.000 ;
    END
  END last_addr[2]
  PIN last_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 745.920 696.000 746.480 700.000 ;
    END
  END last_addr[3]
  PIN last_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 759.360 696.000 759.920 700.000 ;
    END
  END last_addr[4]
  PIN last_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 772.800 696.000 773.360 700.000 ;
    END
  END last_addr[5]
  PIN last_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 786.240 696.000 786.800 700.000 ;
    END
  END last_addr[6]
  PIN last_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 799.680 696.000 800.240 700.000 ;
    END
  END last_addr[7]
  PIN last_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 813.120 696.000 813.680 700.000 ;
    END
  END last_addr[8]
  PIN last_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 826.560 696.000 827.120 700.000 ;
    END
  END last_addr[9]
  PIN le_hi_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 692.160 696.000 692.720 700.000 ;
    END
  END le_hi_act
  PIN le_lo_act
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 678.720 696.000 679.280 700.000 ;
    END
  END le_lo_act
  PIN ram_bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 624.960 4.000 625.520 ;
    END
  END ram_bus_in[0]
  PIN ram_bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 631.680 4.000 632.240 ;
    END
  END ram_bus_in[1]
  PIN ram_bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 638.400 4.000 638.960 ;
    END
  END ram_bus_in[2]
  PIN ram_bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 645.120 4.000 645.680 ;
    END
  END ram_bus_in[3]
  PIN ram_bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 651.840 4.000 652.400 ;
    END
  END ram_bus_in[4]
  PIN ram_bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 658.560 4.000 659.120 ;
    END
  END ram_bus_in[5]
  PIN ram_bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 665.280 4.000 665.840 ;
    END
  END ram_bus_in[6]
  PIN ram_bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.741000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 672.000 4.000 672.560 ;
    END
  END ram_bus_in[7]
  PIN ram_enabled
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 678.720 4.000 679.280 ;
    END
  END ram_enabled
  PIN requested_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 561.120 1050.000 561.680 ;
    END
  END requested_addr[0]
  PIN requested_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 628.320 1050.000 628.880 ;
    END
  END requested_addr[10]
  PIN requested_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 635.040 1050.000 635.600 ;
    END
  END requested_addr[11]
  PIN requested_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 641.760 1050.000 642.320 ;
    END
  END requested_addr[12]
  PIN requested_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 648.480 1050.000 649.040 ;
    END
  END requested_addr[13]
  PIN requested_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 655.200 1050.000 655.760 ;
    END
  END requested_addr[14]
  PIN requested_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 661.920 1050.000 662.480 ;
    END
  END requested_addr[15]
  PIN requested_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 567.840 1050.000 568.400 ;
    END
  END requested_addr[1]
  PIN requested_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 574.560 1050.000 575.120 ;
    END
  END requested_addr[2]
  PIN requested_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 581.280 1050.000 581.840 ;
    END
  END requested_addr[3]
  PIN requested_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 588.000 1050.000 588.560 ;
    END
  END requested_addr[4]
  PIN requested_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 594.720 1050.000 595.280 ;
    END
  END requested_addr[5]
  PIN requested_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 601.440 1050.000 602.000 ;
    END
  END requested_addr[6]
  PIN requested_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 608.160 1050.000 608.720 ;
    END
  END requested_addr[7]
  PIN requested_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 614.880 1050.000 615.440 ;
    END
  END requested_addr[8]
  PIN requested_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 621.600 1050.000 622.160 ;
    END
  END requested_addr[9]
  PIN reset_out
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 1046.000 493.920 1050.000 494.480 ;
    END
  END reset_out
  PIN rom_bus_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 571.200 4.000 571.760 ;
    END
  END rom_bus_in[0]
  PIN rom_bus_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.498500 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 577.920 4.000 578.480 ;
    END
  END rom_bus_in[1]
  PIN rom_bus_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 584.640 4.000 585.200 ;
    END
  END rom_bus_in[2]
  PIN rom_bus_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 591.360 4.000 591.920 ;
    END
  END rom_bus_in[3]
  PIN rom_bus_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 598.080 4.000 598.640 ;
    END
  END rom_bus_in[4]
  PIN rom_bus_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 604.800 4.000 605.360 ;
    END
  END rom_bus_in[5]
  PIN rom_bus_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 611.520 4.000 612.080 ;
    END
  END rom_bus_in[6]
  PIN rom_bus_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.726000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 618.240 4.000 618.800 ;
    END
  END rom_bus_in[7]
  PIN rom_bus_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 517.440 4.000 518.000 ;
    END
  END rom_bus_out[0]
  PIN rom_bus_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 524.160 4.000 524.720 ;
    END
  END rom_bus_out[1]
  PIN rom_bus_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 530.880 4.000 531.440 ;
    END
  END rom_bus_out[2]
  PIN rom_bus_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 537.600 4.000 538.160 ;
    END
  END rom_bus_out[3]
  PIN rom_bus_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 544.320 4.000 544.880 ;
    END
  END rom_bus_out[4]
  PIN rom_bus_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 551.040 4.000 551.600 ;
    END
  END rom_bus_out[5]
  PIN rom_bus_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 557.760 4.000 558.320 ;
    END
  END rom_bus_out[6]
  PIN rom_bus_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 564.480 4.000 565.040 ;
    END
  END rom_bus_out[7]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 329.440 15.380 331.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 483.040 15.380 484.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 636.640 15.380 638.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 790.240 15.380 791.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 943.840 15.380 945.440 682.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 252.640 15.380 254.240 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 406.240 15.380 407.840 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 559.840 15.380 561.440 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 713.440 15.380 715.040 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 867.040 15.380 868.640 682.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 1020.640 15.380 1022.240 682.380 ;
    END
  END vss
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.680 0.000 16.240 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.204000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 25.760 0.000 26.320 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 35.840 0.000 36.400 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 76.160 0.000 76.720 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 378.560 0.000 379.120 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 408.800 0.000 409.360 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 439.040 0.000 439.600 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 469.280 0.000 469.840 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 499.520 0.000 500.080 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 529.760 0.000 530.320 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 560.000 0.000 560.560 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 590.240 0.000 590.800 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 620.480 0.000 621.040 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 650.720 0.000 651.280 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 106.400 0.000 106.960 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 680.960 0.000 681.520 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 711.200 0.000 711.760 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 741.440 0.000 742.000 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 771.680 0.000 772.240 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 801.920 0.000 802.480 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 832.160 0.000 832.720 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 862.400 0.000 862.960 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 892.640 0.000 893.200 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 922.880 0.000 923.440 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 953.120 0.000 953.680 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 136.640 0.000 137.200 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 983.360 0.000 983.920 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 1013.600 0.000 1014.160 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 166.880 0.000 167.440 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 197.120 0.000 197.680 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 227.360 0.000 227.920 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 257.600 0.000 258.160 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 287.840 0.000 288.400 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 318.080 0.000 318.640 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER Metal2 ;
        RECT 348.320 0.000 348.880 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 45.920 0.000 46.480 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 86.240 0.000 86.800 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 388.640 0.000 389.200 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 418.880 0.000 419.440 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 449.120 0.000 449.680 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 479.360 0.000 479.920 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 509.600 0.000 510.160 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 539.840 0.000 540.400 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 570.080 0.000 570.640 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 600.320 0.000 600.880 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 630.560 0.000 631.120 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 660.800 0.000 661.360 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 116.480 0.000 117.040 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 691.040 0.000 691.600 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 721.280 0.000 721.840 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 751.520 0.000 752.080 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 781.760 0.000 782.320 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 812.000 0.000 812.560 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 842.240 0.000 842.800 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 872.480 0.000 873.040 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 902.720 0.000 903.280 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 932.960 0.000 933.520 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 963.200 0.000 963.760 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 146.720 0.000 147.280 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 993.440 0.000 994.000 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 1023.680 0.000 1024.240 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 176.960 0.000 177.520 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 207.200 0.000 207.760 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 237.440 0.000 238.000 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 267.680 0.000 268.240 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 297.920 0.000 298.480 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 328.160 0.000 328.720 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 358.400 0.000 358.960 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 96.320 0.000 96.880 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 398.720 0.000 399.280 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 428.960 0.000 429.520 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 459.200 0.000 459.760 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 489.440 0.000 490.000 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 519.680 0.000 520.240 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 549.920 0.000 550.480 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 580.160 0.000 580.720 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 610.400 0.000 610.960 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 640.640 0.000 641.200 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 670.880 0.000 671.440 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 126.560 0.000 127.120 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 701.120 0.000 701.680 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 731.360 0.000 731.920 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 761.600 0.000 762.160 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 791.840 0.000 792.400 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 822.080 0.000 822.640 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 852.320 0.000 852.880 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 882.560 0.000 883.120 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 912.800 0.000 913.360 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 943.040 0.000 943.600 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 973.280 0.000 973.840 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 156.800 0.000 157.360 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1003.520 0.000 1004.080 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 1033.760 0.000 1034.320 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 187.040 0.000 187.600 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 217.280 0.000 217.840 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 247.520 0.000 248.080 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 277.760 0.000 278.320 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 308.000 0.000 308.560 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 338.240 0.000 338.800 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 368.480 0.000 369.040 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 56.000 0.000 56.560 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.396000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal2 ;
        RECT 66.080 0.000 66.640 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 1043.280 682.380 ;
      LAYER Metal2 ;
        RECT 7.580 695.700 19.860 696.500 ;
        RECT 21.020 695.700 33.300 696.500 ;
        RECT 34.460 695.700 46.740 696.500 ;
        RECT 47.900 695.700 60.180 696.500 ;
        RECT 61.340 695.700 73.620 696.500 ;
        RECT 74.780 695.700 87.060 696.500 ;
        RECT 88.220 695.700 100.500 696.500 ;
        RECT 101.660 695.700 113.940 696.500 ;
        RECT 115.100 695.700 127.380 696.500 ;
        RECT 128.540 695.700 140.820 696.500 ;
        RECT 141.980 695.700 154.260 696.500 ;
        RECT 155.420 695.700 167.700 696.500 ;
        RECT 168.860 695.700 181.140 696.500 ;
        RECT 182.300 695.700 194.580 696.500 ;
        RECT 195.740 695.700 208.020 696.500 ;
        RECT 209.180 695.700 221.460 696.500 ;
        RECT 222.620 695.700 234.900 696.500 ;
        RECT 236.060 695.700 248.340 696.500 ;
        RECT 249.500 695.700 261.780 696.500 ;
        RECT 262.940 695.700 275.220 696.500 ;
        RECT 276.380 695.700 288.660 696.500 ;
        RECT 289.820 695.700 302.100 696.500 ;
        RECT 303.260 695.700 315.540 696.500 ;
        RECT 316.700 695.700 328.980 696.500 ;
        RECT 330.140 695.700 342.420 696.500 ;
        RECT 343.580 695.700 355.860 696.500 ;
        RECT 357.020 695.700 369.300 696.500 ;
        RECT 370.460 695.700 382.740 696.500 ;
        RECT 383.900 695.700 396.180 696.500 ;
        RECT 397.340 695.700 409.620 696.500 ;
        RECT 410.780 695.700 423.060 696.500 ;
        RECT 424.220 695.700 436.500 696.500 ;
        RECT 437.660 695.700 449.940 696.500 ;
        RECT 451.100 695.700 463.380 696.500 ;
        RECT 464.540 695.700 476.820 696.500 ;
        RECT 477.980 695.700 490.260 696.500 ;
        RECT 491.420 695.700 503.700 696.500 ;
        RECT 504.860 695.700 517.140 696.500 ;
        RECT 518.300 695.700 530.580 696.500 ;
        RECT 531.740 695.700 544.020 696.500 ;
        RECT 545.180 695.700 557.460 696.500 ;
        RECT 558.620 695.700 570.900 696.500 ;
        RECT 572.060 695.700 584.340 696.500 ;
        RECT 585.500 695.700 597.780 696.500 ;
        RECT 598.940 695.700 611.220 696.500 ;
        RECT 612.380 695.700 624.660 696.500 ;
        RECT 625.820 695.700 638.100 696.500 ;
        RECT 639.260 695.700 651.540 696.500 ;
        RECT 652.700 695.700 664.980 696.500 ;
        RECT 666.140 695.700 678.420 696.500 ;
        RECT 679.580 695.700 691.860 696.500 ;
        RECT 693.020 695.700 705.300 696.500 ;
        RECT 706.460 695.700 718.740 696.500 ;
        RECT 719.900 695.700 732.180 696.500 ;
        RECT 733.340 695.700 745.620 696.500 ;
        RECT 746.780 695.700 759.060 696.500 ;
        RECT 760.220 695.700 772.500 696.500 ;
        RECT 773.660 695.700 785.940 696.500 ;
        RECT 787.100 695.700 799.380 696.500 ;
        RECT 800.540 695.700 812.820 696.500 ;
        RECT 813.980 695.700 826.260 696.500 ;
        RECT 827.420 695.700 839.700 696.500 ;
        RECT 840.860 695.700 853.140 696.500 ;
        RECT 854.300 695.700 866.580 696.500 ;
        RECT 867.740 695.700 880.020 696.500 ;
        RECT 881.180 695.700 893.460 696.500 ;
        RECT 894.620 695.700 906.900 696.500 ;
        RECT 908.060 695.700 920.340 696.500 ;
        RECT 921.500 695.700 933.780 696.500 ;
        RECT 934.940 695.700 947.220 696.500 ;
        RECT 948.380 695.700 960.660 696.500 ;
        RECT 961.820 695.700 974.100 696.500 ;
        RECT 975.260 695.700 987.540 696.500 ;
        RECT 988.700 695.700 1000.980 696.500 ;
        RECT 1002.140 695.700 1014.420 696.500 ;
        RECT 1015.580 695.700 1027.860 696.500 ;
        RECT 1029.020 695.700 1041.300 696.500 ;
        RECT 1042.460 695.700 1043.700 696.500 ;
        RECT 6.860 4.300 1043.700 695.700 ;
        RECT 6.860 3.500 15.380 4.300 ;
        RECT 16.540 3.500 25.460 4.300 ;
        RECT 26.620 3.500 35.540 4.300 ;
        RECT 36.700 3.500 45.620 4.300 ;
        RECT 46.780 3.500 55.700 4.300 ;
        RECT 56.860 3.500 65.780 4.300 ;
        RECT 66.940 3.500 75.860 4.300 ;
        RECT 77.020 3.500 85.940 4.300 ;
        RECT 87.100 3.500 96.020 4.300 ;
        RECT 97.180 3.500 106.100 4.300 ;
        RECT 107.260 3.500 116.180 4.300 ;
        RECT 117.340 3.500 126.260 4.300 ;
        RECT 127.420 3.500 136.340 4.300 ;
        RECT 137.500 3.500 146.420 4.300 ;
        RECT 147.580 3.500 156.500 4.300 ;
        RECT 157.660 3.500 166.580 4.300 ;
        RECT 167.740 3.500 176.660 4.300 ;
        RECT 177.820 3.500 186.740 4.300 ;
        RECT 187.900 3.500 196.820 4.300 ;
        RECT 197.980 3.500 206.900 4.300 ;
        RECT 208.060 3.500 216.980 4.300 ;
        RECT 218.140 3.500 227.060 4.300 ;
        RECT 228.220 3.500 237.140 4.300 ;
        RECT 238.300 3.500 247.220 4.300 ;
        RECT 248.380 3.500 257.300 4.300 ;
        RECT 258.460 3.500 267.380 4.300 ;
        RECT 268.540 3.500 277.460 4.300 ;
        RECT 278.620 3.500 287.540 4.300 ;
        RECT 288.700 3.500 297.620 4.300 ;
        RECT 298.780 3.500 307.700 4.300 ;
        RECT 308.860 3.500 317.780 4.300 ;
        RECT 318.940 3.500 327.860 4.300 ;
        RECT 329.020 3.500 337.940 4.300 ;
        RECT 339.100 3.500 348.020 4.300 ;
        RECT 349.180 3.500 358.100 4.300 ;
        RECT 359.260 3.500 368.180 4.300 ;
        RECT 369.340 3.500 378.260 4.300 ;
        RECT 379.420 3.500 388.340 4.300 ;
        RECT 389.500 3.500 398.420 4.300 ;
        RECT 399.580 3.500 408.500 4.300 ;
        RECT 409.660 3.500 418.580 4.300 ;
        RECT 419.740 3.500 428.660 4.300 ;
        RECT 429.820 3.500 438.740 4.300 ;
        RECT 439.900 3.500 448.820 4.300 ;
        RECT 449.980 3.500 458.900 4.300 ;
        RECT 460.060 3.500 468.980 4.300 ;
        RECT 470.140 3.500 479.060 4.300 ;
        RECT 480.220 3.500 489.140 4.300 ;
        RECT 490.300 3.500 499.220 4.300 ;
        RECT 500.380 3.500 509.300 4.300 ;
        RECT 510.460 3.500 519.380 4.300 ;
        RECT 520.540 3.500 529.460 4.300 ;
        RECT 530.620 3.500 539.540 4.300 ;
        RECT 540.700 3.500 549.620 4.300 ;
        RECT 550.780 3.500 559.700 4.300 ;
        RECT 560.860 3.500 569.780 4.300 ;
        RECT 570.940 3.500 579.860 4.300 ;
        RECT 581.020 3.500 589.940 4.300 ;
        RECT 591.100 3.500 600.020 4.300 ;
        RECT 601.180 3.500 610.100 4.300 ;
        RECT 611.260 3.500 620.180 4.300 ;
        RECT 621.340 3.500 630.260 4.300 ;
        RECT 631.420 3.500 640.340 4.300 ;
        RECT 641.500 3.500 650.420 4.300 ;
        RECT 651.580 3.500 660.500 4.300 ;
        RECT 661.660 3.500 670.580 4.300 ;
        RECT 671.740 3.500 680.660 4.300 ;
        RECT 681.820 3.500 690.740 4.300 ;
        RECT 691.900 3.500 700.820 4.300 ;
        RECT 701.980 3.500 710.900 4.300 ;
        RECT 712.060 3.500 720.980 4.300 ;
        RECT 722.140 3.500 731.060 4.300 ;
        RECT 732.220 3.500 741.140 4.300 ;
        RECT 742.300 3.500 751.220 4.300 ;
        RECT 752.380 3.500 761.300 4.300 ;
        RECT 762.460 3.500 771.380 4.300 ;
        RECT 772.540 3.500 781.460 4.300 ;
        RECT 782.620 3.500 791.540 4.300 ;
        RECT 792.700 3.500 801.620 4.300 ;
        RECT 802.780 3.500 811.700 4.300 ;
        RECT 812.860 3.500 821.780 4.300 ;
        RECT 822.940 3.500 831.860 4.300 ;
        RECT 833.020 3.500 841.940 4.300 ;
        RECT 843.100 3.500 852.020 4.300 ;
        RECT 853.180 3.500 862.100 4.300 ;
        RECT 863.260 3.500 872.180 4.300 ;
        RECT 873.340 3.500 882.260 4.300 ;
        RECT 883.420 3.500 892.340 4.300 ;
        RECT 893.500 3.500 902.420 4.300 ;
        RECT 903.580 3.500 912.500 4.300 ;
        RECT 913.660 3.500 922.580 4.300 ;
        RECT 923.740 3.500 932.660 4.300 ;
        RECT 933.820 3.500 942.740 4.300 ;
        RECT 943.900 3.500 952.820 4.300 ;
        RECT 953.980 3.500 962.900 4.300 ;
        RECT 964.060 3.500 972.980 4.300 ;
        RECT 974.140 3.500 983.060 4.300 ;
        RECT 984.220 3.500 993.140 4.300 ;
        RECT 994.300 3.500 1003.220 4.300 ;
        RECT 1004.380 3.500 1013.300 4.300 ;
        RECT 1014.460 3.500 1023.380 4.300 ;
        RECT 1024.540 3.500 1033.460 4.300 ;
        RECT 1034.620 3.500 1043.700 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 679.580 1046.500 684.740 ;
        RECT 4.300 678.420 1046.500 679.580 ;
        RECT 4.000 672.860 1046.500 678.420 ;
        RECT 4.300 671.700 1046.500 672.860 ;
        RECT 4.000 666.140 1046.500 671.700 ;
        RECT 4.300 664.980 1046.500 666.140 ;
        RECT 4.000 662.780 1046.500 664.980 ;
        RECT 4.000 661.620 1045.700 662.780 ;
        RECT 4.000 659.420 1046.500 661.620 ;
        RECT 4.300 658.260 1046.500 659.420 ;
        RECT 4.000 656.060 1046.500 658.260 ;
        RECT 4.000 654.900 1045.700 656.060 ;
        RECT 4.000 652.700 1046.500 654.900 ;
        RECT 4.300 651.540 1046.500 652.700 ;
        RECT 4.000 649.340 1046.500 651.540 ;
        RECT 4.000 648.180 1045.700 649.340 ;
        RECT 4.000 645.980 1046.500 648.180 ;
        RECT 4.300 644.820 1046.500 645.980 ;
        RECT 4.000 642.620 1046.500 644.820 ;
        RECT 4.000 641.460 1045.700 642.620 ;
        RECT 4.000 639.260 1046.500 641.460 ;
        RECT 4.300 638.100 1046.500 639.260 ;
        RECT 4.000 635.900 1046.500 638.100 ;
        RECT 4.000 634.740 1045.700 635.900 ;
        RECT 4.000 632.540 1046.500 634.740 ;
        RECT 4.300 631.380 1046.500 632.540 ;
        RECT 4.000 629.180 1046.500 631.380 ;
        RECT 4.000 628.020 1045.700 629.180 ;
        RECT 4.000 625.820 1046.500 628.020 ;
        RECT 4.300 624.660 1046.500 625.820 ;
        RECT 4.000 622.460 1046.500 624.660 ;
        RECT 4.000 621.300 1045.700 622.460 ;
        RECT 4.000 619.100 1046.500 621.300 ;
        RECT 4.300 617.940 1046.500 619.100 ;
        RECT 4.000 615.740 1046.500 617.940 ;
        RECT 4.000 614.580 1045.700 615.740 ;
        RECT 4.000 612.380 1046.500 614.580 ;
        RECT 4.300 611.220 1046.500 612.380 ;
        RECT 4.000 609.020 1046.500 611.220 ;
        RECT 4.000 607.860 1045.700 609.020 ;
        RECT 4.000 605.660 1046.500 607.860 ;
        RECT 4.300 604.500 1046.500 605.660 ;
        RECT 4.000 602.300 1046.500 604.500 ;
        RECT 4.000 601.140 1045.700 602.300 ;
        RECT 4.000 598.940 1046.500 601.140 ;
        RECT 4.300 597.780 1046.500 598.940 ;
        RECT 4.000 595.580 1046.500 597.780 ;
        RECT 4.000 594.420 1045.700 595.580 ;
        RECT 4.000 592.220 1046.500 594.420 ;
        RECT 4.300 591.060 1046.500 592.220 ;
        RECT 4.000 588.860 1046.500 591.060 ;
        RECT 4.000 587.700 1045.700 588.860 ;
        RECT 4.000 585.500 1046.500 587.700 ;
        RECT 4.300 584.340 1046.500 585.500 ;
        RECT 4.000 582.140 1046.500 584.340 ;
        RECT 4.000 580.980 1045.700 582.140 ;
        RECT 4.000 578.780 1046.500 580.980 ;
        RECT 4.300 577.620 1046.500 578.780 ;
        RECT 4.000 575.420 1046.500 577.620 ;
        RECT 4.000 574.260 1045.700 575.420 ;
        RECT 4.000 572.060 1046.500 574.260 ;
        RECT 4.300 570.900 1046.500 572.060 ;
        RECT 4.000 568.700 1046.500 570.900 ;
        RECT 4.000 567.540 1045.700 568.700 ;
        RECT 4.000 565.340 1046.500 567.540 ;
        RECT 4.300 564.180 1046.500 565.340 ;
        RECT 4.000 561.980 1046.500 564.180 ;
        RECT 4.000 560.820 1045.700 561.980 ;
        RECT 4.000 558.620 1046.500 560.820 ;
        RECT 4.300 557.460 1046.500 558.620 ;
        RECT 4.000 555.260 1046.500 557.460 ;
        RECT 4.000 554.100 1045.700 555.260 ;
        RECT 4.000 551.900 1046.500 554.100 ;
        RECT 4.300 550.740 1046.500 551.900 ;
        RECT 4.000 548.540 1046.500 550.740 ;
        RECT 4.000 547.380 1045.700 548.540 ;
        RECT 4.000 545.180 1046.500 547.380 ;
        RECT 4.300 544.020 1046.500 545.180 ;
        RECT 4.000 541.820 1046.500 544.020 ;
        RECT 4.000 540.660 1045.700 541.820 ;
        RECT 4.000 538.460 1046.500 540.660 ;
        RECT 4.300 537.300 1046.500 538.460 ;
        RECT 4.000 535.100 1046.500 537.300 ;
        RECT 4.000 533.940 1045.700 535.100 ;
        RECT 4.000 531.740 1046.500 533.940 ;
        RECT 4.300 530.580 1046.500 531.740 ;
        RECT 4.000 528.380 1046.500 530.580 ;
        RECT 4.000 527.220 1045.700 528.380 ;
        RECT 4.000 525.020 1046.500 527.220 ;
        RECT 4.300 523.860 1046.500 525.020 ;
        RECT 4.000 521.660 1046.500 523.860 ;
        RECT 4.000 520.500 1045.700 521.660 ;
        RECT 4.000 518.300 1046.500 520.500 ;
        RECT 4.300 517.140 1046.500 518.300 ;
        RECT 4.000 514.940 1046.500 517.140 ;
        RECT 4.000 513.780 1045.700 514.940 ;
        RECT 4.000 511.580 1046.500 513.780 ;
        RECT 4.300 510.420 1046.500 511.580 ;
        RECT 4.000 508.220 1046.500 510.420 ;
        RECT 4.000 507.060 1045.700 508.220 ;
        RECT 4.000 504.860 1046.500 507.060 ;
        RECT 4.300 503.700 1046.500 504.860 ;
        RECT 4.000 501.500 1046.500 503.700 ;
        RECT 4.000 500.340 1045.700 501.500 ;
        RECT 4.000 498.140 1046.500 500.340 ;
        RECT 4.300 496.980 1046.500 498.140 ;
        RECT 4.000 494.780 1046.500 496.980 ;
        RECT 4.000 493.620 1045.700 494.780 ;
        RECT 4.000 491.420 1046.500 493.620 ;
        RECT 4.300 490.260 1046.500 491.420 ;
        RECT 4.000 488.060 1046.500 490.260 ;
        RECT 4.000 486.900 1045.700 488.060 ;
        RECT 4.000 484.700 1046.500 486.900 ;
        RECT 4.300 483.540 1046.500 484.700 ;
        RECT 4.000 481.340 1046.500 483.540 ;
        RECT 4.000 480.180 1045.700 481.340 ;
        RECT 4.000 477.980 1046.500 480.180 ;
        RECT 4.300 476.820 1046.500 477.980 ;
        RECT 4.000 474.620 1046.500 476.820 ;
        RECT 4.000 473.460 1045.700 474.620 ;
        RECT 4.000 471.260 1046.500 473.460 ;
        RECT 4.300 470.100 1046.500 471.260 ;
        RECT 4.000 467.900 1046.500 470.100 ;
        RECT 4.000 466.740 1045.700 467.900 ;
        RECT 4.000 464.540 1046.500 466.740 ;
        RECT 4.300 463.380 1046.500 464.540 ;
        RECT 4.000 461.180 1046.500 463.380 ;
        RECT 4.000 460.020 1045.700 461.180 ;
        RECT 4.000 457.820 1046.500 460.020 ;
        RECT 4.300 456.660 1046.500 457.820 ;
        RECT 4.000 454.460 1046.500 456.660 ;
        RECT 4.000 453.300 1045.700 454.460 ;
        RECT 4.000 451.100 1046.500 453.300 ;
        RECT 4.300 449.940 1046.500 451.100 ;
        RECT 4.000 447.740 1046.500 449.940 ;
        RECT 4.000 446.580 1045.700 447.740 ;
        RECT 4.000 444.380 1046.500 446.580 ;
        RECT 4.300 443.220 1046.500 444.380 ;
        RECT 4.000 441.020 1046.500 443.220 ;
        RECT 4.000 439.860 1045.700 441.020 ;
        RECT 4.000 437.660 1046.500 439.860 ;
        RECT 4.300 436.500 1046.500 437.660 ;
        RECT 4.000 434.300 1046.500 436.500 ;
        RECT 4.000 433.140 1045.700 434.300 ;
        RECT 4.000 430.940 1046.500 433.140 ;
        RECT 4.300 429.780 1046.500 430.940 ;
        RECT 4.000 427.580 1046.500 429.780 ;
        RECT 4.000 426.420 1045.700 427.580 ;
        RECT 4.000 424.220 1046.500 426.420 ;
        RECT 4.300 423.060 1046.500 424.220 ;
        RECT 4.000 420.860 1046.500 423.060 ;
        RECT 4.000 419.700 1045.700 420.860 ;
        RECT 4.000 417.500 1046.500 419.700 ;
        RECT 4.300 416.340 1046.500 417.500 ;
        RECT 4.000 414.140 1046.500 416.340 ;
        RECT 4.000 412.980 1045.700 414.140 ;
        RECT 4.000 410.780 1046.500 412.980 ;
        RECT 4.300 409.620 1046.500 410.780 ;
        RECT 4.000 407.420 1046.500 409.620 ;
        RECT 4.000 406.260 1045.700 407.420 ;
        RECT 4.000 404.060 1046.500 406.260 ;
        RECT 4.300 402.900 1046.500 404.060 ;
        RECT 4.000 400.700 1046.500 402.900 ;
        RECT 4.000 399.540 1045.700 400.700 ;
        RECT 4.000 397.340 1046.500 399.540 ;
        RECT 4.300 396.180 1046.500 397.340 ;
        RECT 4.000 393.980 1046.500 396.180 ;
        RECT 4.000 392.820 1045.700 393.980 ;
        RECT 4.000 390.620 1046.500 392.820 ;
        RECT 4.300 389.460 1046.500 390.620 ;
        RECT 4.000 387.260 1046.500 389.460 ;
        RECT 4.000 386.100 1045.700 387.260 ;
        RECT 4.000 383.900 1046.500 386.100 ;
        RECT 4.300 382.740 1046.500 383.900 ;
        RECT 4.000 380.540 1046.500 382.740 ;
        RECT 4.000 379.380 1045.700 380.540 ;
        RECT 4.000 377.180 1046.500 379.380 ;
        RECT 4.300 376.020 1046.500 377.180 ;
        RECT 4.000 373.820 1046.500 376.020 ;
        RECT 4.000 372.660 1045.700 373.820 ;
        RECT 4.000 370.460 1046.500 372.660 ;
        RECT 4.300 369.300 1046.500 370.460 ;
        RECT 4.000 367.100 1046.500 369.300 ;
        RECT 4.000 365.940 1045.700 367.100 ;
        RECT 4.000 363.740 1046.500 365.940 ;
        RECT 4.300 362.580 1046.500 363.740 ;
        RECT 4.000 360.380 1046.500 362.580 ;
        RECT 4.000 359.220 1045.700 360.380 ;
        RECT 4.000 357.020 1046.500 359.220 ;
        RECT 4.300 355.860 1046.500 357.020 ;
        RECT 4.000 353.660 1046.500 355.860 ;
        RECT 4.000 352.500 1045.700 353.660 ;
        RECT 4.000 350.300 1046.500 352.500 ;
        RECT 4.300 349.140 1046.500 350.300 ;
        RECT 4.000 346.940 1046.500 349.140 ;
        RECT 4.000 345.780 1045.700 346.940 ;
        RECT 4.000 343.580 1046.500 345.780 ;
        RECT 4.300 342.420 1046.500 343.580 ;
        RECT 4.000 340.220 1046.500 342.420 ;
        RECT 4.000 339.060 1045.700 340.220 ;
        RECT 4.000 336.860 1046.500 339.060 ;
        RECT 4.300 335.700 1046.500 336.860 ;
        RECT 4.000 333.500 1046.500 335.700 ;
        RECT 4.000 332.340 1045.700 333.500 ;
        RECT 4.000 330.140 1046.500 332.340 ;
        RECT 4.300 328.980 1046.500 330.140 ;
        RECT 4.000 326.780 1046.500 328.980 ;
        RECT 4.000 325.620 1045.700 326.780 ;
        RECT 4.000 323.420 1046.500 325.620 ;
        RECT 4.300 322.260 1046.500 323.420 ;
        RECT 4.000 320.060 1046.500 322.260 ;
        RECT 4.000 318.900 1045.700 320.060 ;
        RECT 4.000 316.700 1046.500 318.900 ;
        RECT 4.300 315.540 1046.500 316.700 ;
        RECT 4.000 313.340 1046.500 315.540 ;
        RECT 4.000 312.180 1045.700 313.340 ;
        RECT 4.000 309.980 1046.500 312.180 ;
        RECT 4.300 308.820 1046.500 309.980 ;
        RECT 4.000 306.620 1046.500 308.820 ;
        RECT 4.000 305.460 1045.700 306.620 ;
        RECT 4.000 303.260 1046.500 305.460 ;
        RECT 4.300 302.100 1046.500 303.260 ;
        RECT 4.000 299.900 1046.500 302.100 ;
        RECT 4.000 298.740 1045.700 299.900 ;
        RECT 4.000 296.540 1046.500 298.740 ;
        RECT 4.300 295.380 1046.500 296.540 ;
        RECT 4.000 293.180 1046.500 295.380 ;
        RECT 4.000 292.020 1045.700 293.180 ;
        RECT 4.000 289.820 1046.500 292.020 ;
        RECT 4.300 288.660 1046.500 289.820 ;
        RECT 4.000 286.460 1046.500 288.660 ;
        RECT 4.000 285.300 1045.700 286.460 ;
        RECT 4.000 283.100 1046.500 285.300 ;
        RECT 4.300 281.940 1046.500 283.100 ;
        RECT 4.000 279.740 1046.500 281.940 ;
        RECT 4.000 278.580 1045.700 279.740 ;
        RECT 4.000 276.380 1046.500 278.580 ;
        RECT 4.300 275.220 1046.500 276.380 ;
        RECT 4.000 273.020 1046.500 275.220 ;
        RECT 4.000 271.860 1045.700 273.020 ;
        RECT 4.000 269.660 1046.500 271.860 ;
        RECT 4.300 268.500 1046.500 269.660 ;
        RECT 4.000 266.300 1046.500 268.500 ;
        RECT 4.000 265.140 1045.700 266.300 ;
        RECT 4.000 262.940 1046.500 265.140 ;
        RECT 4.300 261.780 1046.500 262.940 ;
        RECT 4.000 259.580 1046.500 261.780 ;
        RECT 4.000 258.420 1045.700 259.580 ;
        RECT 4.000 256.220 1046.500 258.420 ;
        RECT 4.300 255.060 1046.500 256.220 ;
        RECT 4.000 252.860 1046.500 255.060 ;
        RECT 4.000 251.700 1045.700 252.860 ;
        RECT 4.000 249.500 1046.500 251.700 ;
        RECT 4.300 248.340 1046.500 249.500 ;
        RECT 4.000 246.140 1046.500 248.340 ;
        RECT 4.000 244.980 1045.700 246.140 ;
        RECT 4.000 242.780 1046.500 244.980 ;
        RECT 4.300 241.620 1046.500 242.780 ;
        RECT 4.000 239.420 1046.500 241.620 ;
        RECT 4.000 238.260 1045.700 239.420 ;
        RECT 4.000 236.060 1046.500 238.260 ;
        RECT 4.300 234.900 1046.500 236.060 ;
        RECT 4.000 232.700 1046.500 234.900 ;
        RECT 4.000 231.540 1045.700 232.700 ;
        RECT 4.000 229.340 1046.500 231.540 ;
        RECT 4.300 228.180 1046.500 229.340 ;
        RECT 4.000 225.980 1046.500 228.180 ;
        RECT 4.000 224.820 1045.700 225.980 ;
        RECT 4.000 222.620 1046.500 224.820 ;
        RECT 4.300 221.460 1046.500 222.620 ;
        RECT 4.000 219.260 1046.500 221.460 ;
        RECT 4.000 218.100 1045.700 219.260 ;
        RECT 4.000 215.900 1046.500 218.100 ;
        RECT 4.300 214.740 1046.500 215.900 ;
        RECT 4.000 212.540 1046.500 214.740 ;
        RECT 4.000 211.380 1045.700 212.540 ;
        RECT 4.000 209.180 1046.500 211.380 ;
        RECT 4.300 208.020 1046.500 209.180 ;
        RECT 4.000 205.820 1046.500 208.020 ;
        RECT 4.000 204.660 1045.700 205.820 ;
        RECT 4.000 202.460 1046.500 204.660 ;
        RECT 4.300 201.300 1046.500 202.460 ;
        RECT 4.000 199.100 1046.500 201.300 ;
        RECT 4.000 197.940 1045.700 199.100 ;
        RECT 4.000 195.740 1046.500 197.940 ;
        RECT 4.300 194.580 1046.500 195.740 ;
        RECT 4.000 192.380 1046.500 194.580 ;
        RECT 4.000 191.220 1045.700 192.380 ;
        RECT 4.000 189.020 1046.500 191.220 ;
        RECT 4.300 187.860 1046.500 189.020 ;
        RECT 4.000 185.660 1046.500 187.860 ;
        RECT 4.000 184.500 1045.700 185.660 ;
        RECT 4.000 182.300 1046.500 184.500 ;
        RECT 4.300 181.140 1046.500 182.300 ;
        RECT 4.000 178.940 1046.500 181.140 ;
        RECT 4.000 177.780 1045.700 178.940 ;
        RECT 4.000 175.580 1046.500 177.780 ;
        RECT 4.300 174.420 1046.500 175.580 ;
        RECT 4.000 172.220 1046.500 174.420 ;
        RECT 4.000 171.060 1045.700 172.220 ;
        RECT 4.000 168.860 1046.500 171.060 ;
        RECT 4.300 167.700 1046.500 168.860 ;
        RECT 4.000 165.500 1046.500 167.700 ;
        RECT 4.000 164.340 1045.700 165.500 ;
        RECT 4.000 162.140 1046.500 164.340 ;
        RECT 4.300 160.980 1046.500 162.140 ;
        RECT 4.000 158.780 1046.500 160.980 ;
        RECT 4.000 157.620 1045.700 158.780 ;
        RECT 4.000 155.420 1046.500 157.620 ;
        RECT 4.300 154.260 1046.500 155.420 ;
        RECT 4.000 152.060 1046.500 154.260 ;
        RECT 4.000 150.900 1045.700 152.060 ;
        RECT 4.000 148.700 1046.500 150.900 ;
        RECT 4.300 147.540 1046.500 148.700 ;
        RECT 4.000 145.340 1046.500 147.540 ;
        RECT 4.000 144.180 1045.700 145.340 ;
        RECT 4.000 141.980 1046.500 144.180 ;
        RECT 4.300 140.820 1046.500 141.980 ;
        RECT 4.000 138.620 1046.500 140.820 ;
        RECT 4.000 137.460 1045.700 138.620 ;
        RECT 4.000 135.260 1046.500 137.460 ;
        RECT 4.300 134.100 1046.500 135.260 ;
        RECT 4.000 131.900 1046.500 134.100 ;
        RECT 4.000 130.740 1045.700 131.900 ;
        RECT 4.000 128.540 1046.500 130.740 ;
        RECT 4.300 127.380 1046.500 128.540 ;
        RECT 4.000 125.180 1046.500 127.380 ;
        RECT 4.000 124.020 1045.700 125.180 ;
        RECT 4.000 121.820 1046.500 124.020 ;
        RECT 4.300 120.660 1046.500 121.820 ;
        RECT 4.000 118.460 1046.500 120.660 ;
        RECT 4.000 117.300 1045.700 118.460 ;
        RECT 4.000 115.100 1046.500 117.300 ;
        RECT 4.300 113.940 1046.500 115.100 ;
        RECT 4.000 111.740 1046.500 113.940 ;
        RECT 4.000 110.580 1045.700 111.740 ;
        RECT 4.000 108.380 1046.500 110.580 ;
        RECT 4.300 107.220 1046.500 108.380 ;
        RECT 4.000 105.020 1046.500 107.220 ;
        RECT 4.000 103.860 1045.700 105.020 ;
        RECT 4.000 101.660 1046.500 103.860 ;
        RECT 4.300 100.500 1046.500 101.660 ;
        RECT 4.000 98.300 1046.500 100.500 ;
        RECT 4.000 97.140 1045.700 98.300 ;
        RECT 4.000 94.940 1046.500 97.140 ;
        RECT 4.300 93.780 1046.500 94.940 ;
        RECT 4.000 91.580 1046.500 93.780 ;
        RECT 4.000 90.420 1045.700 91.580 ;
        RECT 4.000 88.220 1046.500 90.420 ;
        RECT 4.300 87.060 1046.500 88.220 ;
        RECT 4.000 84.860 1046.500 87.060 ;
        RECT 4.000 83.700 1045.700 84.860 ;
        RECT 4.000 81.500 1046.500 83.700 ;
        RECT 4.300 80.340 1046.500 81.500 ;
        RECT 4.000 78.140 1046.500 80.340 ;
        RECT 4.000 76.980 1045.700 78.140 ;
        RECT 4.000 74.780 1046.500 76.980 ;
        RECT 4.300 73.620 1046.500 74.780 ;
        RECT 4.000 71.420 1046.500 73.620 ;
        RECT 4.000 70.260 1045.700 71.420 ;
        RECT 4.000 68.060 1046.500 70.260 ;
        RECT 4.300 66.900 1046.500 68.060 ;
        RECT 4.000 64.700 1046.500 66.900 ;
        RECT 4.000 63.540 1045.700 64.700 ;
        RECT 4.000 61.340 1046.500 63.540 ;
        RECT 4.300 60.180 1046.500 61.340 ;
        RECT 4.000 57.980 1046.500 60.180 ;
        RECT 4.000 56.820 1045.700 57.980 ;
        RECT 4.000 54.620 1046.500 56.820 ;
        RECT 4.300 53.460 1046.500 54.620 ;
        RECT 4.000 51.260 1046.500 53.460 ;
        RECT 4.000 50.100 1045.700 51.260 ;
        RECT 4.000 47.900 1046.500 50.100 ;
        RECT 4.300 46.740 1046.500 47.900 ;
        RECT 4.000 44.540 1046.500 46.740 ;
        RECT 4.000 43.380 1045.700 44.540 ;
        RECT 4.000 41.180 1046.500 43.380 ;
        RECT 4.300 40.020 1046.500 41.180 ;
        RECT 4.000 37.820 1046.500 40.020 ;
        RECT 4.000 36.660 1045.700 37.820 ;
        RECT 4.000 34.460 1046.500 36.660 ;
        RECT 4.300 33.300 1046.500 34.460 ;
        RECT 4.000 27.740 1046.500 33.300 ;
        RECT 4.300 26.580 1046.500 27.740 ;
        RECT 4.000 21.020 1046.500 26.580 ;
        RECT 4.300 19.860 1046.500 21.020 ;
        RECT 4.000 14.140 1046.500 19.860 ;
      LAYER Metal4 ;
        RECT 130.620 60.010 175.540 665.750 ;
        RECT 177.740 60.010 252.340 665.750 ;
        RECT 254.540 60.010 329.140 665.750 ;
        RECT 331.340 60.010 405.940 665.750 ;
        RECT 408.140 60.010 482.740 665.750 ;
        RECT 484.940 60.010 559.540 665.750 ;
        RECT 561.740 60.010 636.340 665.750 ;
        RECT 638.540 60.010 713.140 665.750 ;
        RECT 715.340 60.010 789.940 665.750 ;
        RECT 792.140 60.010 866.740 665.750 ;
        RECT 868.940 60.010 943.540 665.750 ;
        RECT 945.740 60.010 998.900 665.750 ;
  END
END wrapped_as2650
END LIBRARY

