magic
tech gf180mcuD
magscale 1 10
timestamp 1701963850
<< metal2 >>
rect 3744 98504 3856 99176
rect 3724 98376 3856 98504
rect 4444 98504 4556 99176
rect 5344 98504 5456 99176
rect 4444 98376 4564 98504
rect 5344 98376 5460 98504
rect 13444 98376 13556 99176
rect 14144 98504 14256 99176
rect 14140 98376 14256 98504
rect 14544 98376 14656 99176
rect 14994 98376 15106 99176
rect 15444 98376 15556 99176
rect 16044 98376 16156 99176
rect 24244 98504 24356 99176
rect 24220 98376 24356 98504
rect 25044 98504 25156 99176
rect 25044 98376 25172 98504
rect 25744 98376 25856 99176
rect 30944 98504 31056 99176
rect 30940 98376 31056 98504
rect 31944 98376 32056 99176
rect 32744 98504 32856 99176
rect 32732 98376 32856 98504
rect 33344 98504 33456 99176
rect 33344 98376 33460 98504
rect 36844 98376 36956 99176
rect 46568 98376 46680 99176
rect 52944 98504 53056 99176
rect 52944 98376 53060 98504
rect 54644 98376 54756 99176
rect 56344 98376 56456 99176
rect 57444 98376 57556 99176
rect 58144 98376 58256 99176
rect 59244 98376 59356 99176
rect 63344 98504 63456 99176
rect 63344 98376 63476 98504
rect 63744 98376 63856 99176
rect 64944 98376 65056 99176
rect 73044 98376 73156 99176
rect 73744 98504 73856 99176
rect 73724 98376 73856 98504
rect 74144 98376 74256 99176
rect 74544 98504 74656 99176
rect 74544 98376 74676 98504
rect 74944 98376 75056 99176
rect 75644 98504 75756 99176
rect 75628 98376 75756 98504
rect 83844 98504 83956 99176
rect 83844 98376 83972 98504
rect 84644 98376 84756 99176
rect 85344 98376 85456 99176
rect 3724 98196 3780 98376
rect 3724 98140 3836 98196
rect 3780 97944 3836 98140
rect 4508 97944 4564 98376
rect 5404 97944 5460 98376
rect 13468 97944 13524 98376
rect 14140 97944 14196 98376
rect 14588 97944 14644 98376
rect 15036 97944 15092 98376
rect 15484 97944 15540 98376
rect 16044 97944 16100 98376
rect 24220 97944 24276 98376
rect 25116 97944 25172 98376
rect 25788 97944 25844 98376
rect 30940 97944 30996 98376
rect 31948 98196 32004 98376
rect 31948 98140 32060 98196
rect 32004 97944 32060 98140
rect 32732 97944 32788 98376
rect 33404 97944 33460 98376
rect 36876 97944 36932 98376
rect 46620 97944 46676 98376
rect 53004 97944 53060 98376
rect 54684 97944 54740 98376
rect 56364 97944 56420 98376
rect 57484 97944 57540 98376
rect 58156 97944 58212 98376
rect 59276 97944 59332 98376
rect 63420 97944 63476 98376
rect 63756 97944 63812 98376
rect 64988 97944 65044 98376
rect 73052 97944 73108 98376
rect 73724 97944 73780 98376
rect 74172 97944 74228 98376
rect 74620 97944 74676 98376
rect 74956 97944 75012 98376
rect 75628 97944 75684 98376
rect 83916 97944 83972 98376
rect 84700 97944 84756 98376
rect 85372 97944 85428 98376
<< metal3 >>
rect 1844 95425 2014 95474
rect 1844 95369 1901 95425
rect 1957 95369 2014 95425
rect 1844 95301 2014 95369
rect 1844 95245 1901 95301
rect 1957 95245 2014 95301
rect 1844 95177 2014 95245
rect 1844 95121 1901 95177
rect 1957 95121 2014 95177
rect 1844 95053 2014 95121
rect 1844 94997 1901 95053
rect 1957 94997 2014 95053
rect 1844 94929 2014 94997
rect 1844 94873 1901 94929
rect 1957 94873 2014 94929
rect 1844 94805 2014 94873
rect 1844 94749 1901 94805
rect 1957 94749 2014 94805
rect 1844 94681 2014 94749
rect 1844 94625 1901 94681
rect 1957 94625 2014 94681
rect 1844 94557 2014 94625
rect 1844 94501 1901 94557
rect 1957 94501 2014 94557
rect 1844 94433 2014 94501
rect 1844 94377 1901 94433
rect 1957 94377 2014 94433
rect 1844 94309 2014 94377
rect 1844 94253 1901 94309
rect 1957 94253 2014 94309
rect 1844 94204 2014 94253
rect 86526 95425 86630 95474
rect 86526 95369 86550 95425
rect 86606 95369 86630 95425
rect 86526 95301 86630 95369
rect 86526 95245 86550 95301
rect 86606 95245 86630 95301
rect 86526 95177 86630 95245
rect 86526 95121 86550 95177
rect 86606 95121 86630 95177
rect 86526 95053 86630 95121
rect 86526 94997 86550 95053
rect 86606 94997 86630 95053
rect 86526 94929 86630 94997
rect 86526 94873 86550 94929
rect 86606 94873 86630 94929
rect 86526 94805 86630 94873
rect 86526 94749 86550 94805
rect 86606 94749 86630 94805
rect 86526 94681 86630 94749
rect 86526 94625 86550 94681
rect 86606 94625 86630 94681
rect 86526 94557 86630 94625
rect 86526 94501 86550 94557
rect 86606 94501 86630 94557
rect 86526 94433 86630 94501
rect 86526 94377 86550 94433
rect 86606 94377 86630 94433
rect 86526 94309 86630 94377
rect 86526 94253 86550 94309
rect 86606 94253 86630 94309
rect 86526 94204 86630 94253
rect 86650 95425 87126 95474
rect 86650 95369 86674 95425
rect 86730 95369 86798 95425
rect 86854 95369 86922 95425
rect 86978 95369 87046 95425
rect 87102 95369 87126 95425
rect 86650 95301 87126 95369
rect 86650 95245 86674 95301
rect 86730 95245 86798 95301
rect 86854 95245 86922 95301
rect 86978 95245 87046 95301
rect 87102 95245 87126 95301
rect 86650 95177 87126 95245
rect 86650 95121 86674 95177
rect 86730 95121 86798 95177
rect 86854 95121 86922 95177
rect 86978 95121 87046 95177
rect 87102 95121 87126 95177
rect 86650 95053 87126 95121
rect 86650 94997 86674 95053
rect 86730 94997 86798 95053
rect 86854 94997 86922 95053
rect 86978 94997 87046 95053
rect 87102 94997 87126 95053
rect 86650 94929 87126 94997
rect 86650 94873 86674 94929
rect 86730 94873 86798 94929
rect 86854 94873 86922 94929
rect 86978 94873 87046 94929
rect 87102 94873 87126 94929
rect 86650 94805 87126 94873
rect 86650 94749 86674 94805
rect 86730 94749 86798 94805
rect 86854 94749 86922 94805
rect 86978 94749 87046 94805
rect 87102 94749 87126 94805
rect 86650 94681 87126 94749
rect 86650 94625 86674 94681
rect 86730 94625 86798 94681
rect 86854 94625 86922 94681
rect 86978 94625 87046 94681
rect 87102 94625 87126 94681
rect 86650 94557 87126 94625
rect 86650 94501 86674 94557
rect 86730 94501 86798 94557
rect 86854 94501 86922 94557
rect 86978 94501 87046 94557
rect 87102 94501 87126 94557
rect 86650 94433 87126 94501
rect 86650 94377 86674 94433
rect 86730 94377 86798 94433
rect 86854 94377 86922 94433
rect 86978 94377 87046 94433
rect 87102 94377 87126 94433
rect 86650 94309 87126 94377
rect 86650 94253 86674 94309
rect 86730 94253 86798 94309
rect 86854 94253 86922 94309
rect 86978 94253 87046 94309
rect 87102 94253 87126 94309
rect 86650 94204 87126 94253
rect 86526 92191 86630 92210
rect 86526 92135 86550 92191
rect 86606 92135 86630 92191
rect 86526 92067 86630 92135
rect 86526 92011 86550 92067
rect 86606 92011 86630 92067
rect 86526 91943 86630 92011
rect 86526 91887 86550 91943
rect 86606 91887 86630 91943
rect 86526 91819 86630 91887
rect 86526 91763 86550 91819
rect 86606 91763 86630 91819
rect 86526 91744 86630 91763
rect 86650 92191 87126 92210
rect 86650 92135 86674 92191
rect 86730 92135 86798 92191
rect 86854 92135 86922 92191
rect 86978 92135 87046 92191
rect 87102 92135 87126 92191
rect 86650 92067 87126 92135
rect 86650 92011 86674 92067
rect 86730 92011 86798 92067
rect 86854 92011 86922 92067
rect 86978 92011 87046 92067
rect 87102 92011 87126 92067
rect 86650 91943 87126 92011
rect 86650 91887 86674 91943
rect 86730 91887 86798 91943
rect 86854 91887 86922 91943
rect 86978 91887 87046 91943
rect 87102 91887 87126 91943
rect 86650 91819 87126 91887
rect 86650 91763 86674 91819
rect 86730 91763 86798 91819
rect 86854 91763 86922 91819
rect 86978 91763 87046 91819
rect 87102 91763 87126 91819
rect 86650 91744 87126 91763
rect 86526 91695 86630 91714
rect 86526 91639 86550 91695
rect 86606 91639 86630 91695
rect 86526 91571 86630 91639
rect 86526 91515 86550 91571
rect 86606 91515 86630 91571
rect 86526 91447 86630 91515
rect 86526 91391 86550 91447
rect 86606 91391 86630 91447
rect 86526 91323 86630 91391
rect 86526 91267 86550 91323
rect 86606 91267 86630 91323
rect 86526 91248 86630 91267
rect 86650 91695 87126 91714
rect 86650 91639 86674 91695
rect 86730 91639 86798 91695
rect 86854 91639 86922 91695
rect 86978 91639 87046 91695
rect 87102 91639 87126 91695
rect 86650 91571 87126 91639
rect 86650 91515 86674 91571
rect 86730 91515 86798 91571
rect 86854 91515 86922 91571
rect 86978 91515 87046 91571
rect 87102 91515 87126 91571
rect 86650 91447 87126 91515
rect 86650 91391 86674 91447
rect 86730 91391 86798 91447
rect 86854 91391 86922 91447
rect 86978 91391 87046 91447
rect 87102 91391 87126 91447
rect 86650 91323 87126 91391
rect 86650 91267 86674 91323
rect 86730 91267 86798 91323
rect 86854 91267 86922 91323
rect 86978 91267 87046 91323
rect 87102 91267 87126 91323
rect 86650 91248 87126 91267
rect 86526 91199 86630 91218
rect 86526 91143 86550 91199
rect 86606 91143 86630 91199
rect 86526 91075 86630 91143
rect 86526 91019 86550 91075
rect 86606 91019 86630 91075
rect 86526 90951 86630 91019
rect 1906 90901 2382 90932
rect 1906 90845 1930 90901
rect 1986 90845 2054 90901
rect 2110 90845 2178 90901
rect 2234 90845 2302 90901
rect 2358 90845 2382 90901
rect 1906 90777 2382 90845
rect 1906 90721 1930 90777
rect 1986 90721 2054 90777
rect 2110 90721 2178 90777
rect 2234 90721 2302 90777
rect 2358 90721 2382 90777
rect 86526 90895 86550 90951
rect 86606 90895 86630 90951
rect 86526 90827 86630 90895
rect 86526 90771 86550 90827
rect 86606 90771 86630 90827
rect 86526 90752 86630 90771
rect 86650 91199 87126 91218
rect 86650 91143 86674 91199
rect 86730 91143 86798 91199
rect 86854 91143 86922 91199
rect 86978 91143 87046 91199
rect 87102 91143 87126 91199
rect 86650 91075 87126 91143
rect 86650 91019 86674 91075
rect 86730 91019 86798 91075
rect 86854 91019 86922 91075
rect 86978 91019 87046 91075
rect 87102 91019 87126 91075
rect 86650 90951 87126 91019
rect 86650 90895 86674 90951
rect 86730 90895 86798 90951
rect 86854 90895 86922 90951
rect 86978 90895 87046 90951
rect 87102 90895 87126 90951
rect 86650 90827 87126 90895
rect 86650 90771 86674 90827
rect 86730 90771 86798 90827
rect 86854 90771 86922 90827
rect 86978 90771 87046 90827
rect 87102 90771 87126 90827
rect 86650 90752 87126 90771
rect 1906 90653 2382 90721
rect 1906 90597 1930 90653
rect 1986 90597 2054 90653
rect 2110 90597 2178 90653
rect 2234 90597 2302 90653
rect 2358 90597 2382 90653
rect 1906 90529 2382 90597
rect 1906 90473 1930 90529
rect 1986 90473 2054 90529
rect 2110 90473 2178 90529
rect 2234 90473 2302 90529
rect 2358 90473 2382 90529
rect 1906 90442 2382 90473
rect 86526 90703 86630 90722
rect 86526 90647 86550 90703
rect 86606 90647 86630 90703
rect 86526 90579 86630 90647
rect 86526 90523 86550 90579
rect 86606 90523 86630 90579
rect 86526 90455 86630 90523
rect 86526 90399 86550 90455
rect 86606 90399 86630 90455
rect 86526 90380 86630 90399
rect 86650 90703 87126 90722
rect 86650 90647 86674 90703
rect 86730 90647 86798 90703
rect 86854 90647 86922 90703
rect 86978 90647 87046 90703
rect 87102 90647 87126 90703
rect 86650 90579 87126 90647
rect 86650 90523 86674 90579
rect 86730 90523 86798 90579
rect 86854 90523 86922 90579
rect 86978 90523 87046 90579
rect 87102 90523 87126 90579
rect 86650 90455 87126 90523
rect 86650 90399 86674 90455
rect 86730 90399 86798 90455
rect 86854 90399 86922 90455
rect 86978 90399 87046 90455
rect 87102 90399 87126 90455
rect 86650 90380 87126 90399
rect 85726 89791 85830 89824
rect 85726 89735 85750 89791
rect 85806 89735 85830 89791
rect 85726 89667 85830 89735
rect 85726 89611 85750 89667
rect 85806 89611 85830 89667
rect 85726 89543 85830 89611
rect 85726 89487 85750 89543
rect 85806 89487 85830 89543
rect 85726 89419 85830 89487
rect 85726 89363 85750 89419
rect 85806 89363 85830 89419
rect 85726 89330 85830 89363
rect 85850 89791 86326 89824
rect 85850 89735 85874 89791
rect 85930 89735 85998 89791
rect 86054 89735 86122 89791
rect 86178 89735 86246 89791
rect 86302 89735 86326 89791
rect 85850 89667 86326 89735
rect 85850 89611 85874 89667
rect 85930 89611 85998 89667
rect 86054 89611 86122 89667
rect 86178 89611 86246 89667
rect 86302 89611 86326 89667
rect 85850 89543 86326 89611
rect 85850 89487 85874 89543
rect 85930 89487 85998 89543
rect 86054 89487 86122 89543
rect 86178 89487 86246 89543
rect 86302 89487 86326 89543
rect 85850 89419 86326 89487
rect 85850 89363 85874 89419
rect 85930 89363 85998 89419
rect 86054 89363 86122 89419
rect 86178 89363 86246 89419
rect 86302 89363 86326 89419
rect 85850 89330 86326 89363
rect 85726 89295 85830 89328
rect 85726 89239 85750 89295
rect 85806 89239 85830 89295
rect 85726 89171 85830 89239
rect 85726 89115 85750 89171
rect 85806 89115 85830 89171
rect 85726 89047 85830 89115
rect 85726 88991 85750 89047
rect 85806 88991 85830 89047
rect 85726 88923 85830 88991
rect 85726 88867 85750 88923
rect 85806 88867 85830 88923
rect 85726 88834 85830 88867
rect 85850 89295 86326 89328
rect 85850 89239 85874 89295
rect 85930 89239 85998 89295
rect 86054 89239 86122 89295
rect 86178 89239 86246 89295
rect 86302 89239 86326 89295
rect 85850 89171 86326 89239
rect 85850 89115 85874 89171
rect 85930 89115 85998 89171
rect 86054 89115 86122 89171
rect 86178 89115 86246 89171
rect 86302 89115 86326 89171
rect 85850 89047 86326 89115
rect 85850 88991 85874 89047
rect 85930 88991 85998 89047
rect 86054 88991 86122 89047
rect 86178 88991 86246 89047
rect 86302 88991 86326 89047
rect 85850 88923 86326 88991
rect 85850 88867 85874 88923
rect 85930 88867 85998 88923
rect 86054 88867 86122 88923
rect 86178 88867 86246 88923
rect 86302 88867 86326 88923
rect 85850 88834 86326 88867
rect 85726 88799 85830 88832
rect 85726 88743 85750 88799
rect 85806 88743 85830 88799
rect 85726 88675 85830 88743
rect 85726 88619 85750 88675
rect 85806 88619 85830 88675
rect 85726 88551 85830 88619
rect 85726 88495 85750 88551
rect 85806 88495 85830 88551
rect 85726 88462 85830 88495
rect 85850 88799 86326 88832
rect 85850 88743 85874 88799
rect 85930 88743 85998 88799
rect 86054 88743 86122 88799
rect 86178 88743 86246 88799
rect 86302 88743 86326 88799
rect 85850 88675 86326 88743
rect 85850 88619 85874 88675
rect 85930 88619 85998 88675
rect 86054 88619 86122 88675
rect 86178 88619 86246 88675
rect 86302 88619 86326 88675
rect 85850 88551 86326 88619
rect 85850 88495 85874 88551
rect 85930 88495 85998 88551
rect 86054 88495 86122 88551
rect 86178 88495 86246 88551
rect 86302 88495 86326 88551
rect 85850 88462 86326 88495
rect 1044 85889 1148 85940
rect 1044 85833 1068 85889
rect 1124 85833 1148 85889
rect 1044 85765 1148 85833
rect 1044 85709 1068 85765
rect 1124 85709 1148 85765
rect 1044 85641 1148 85709
rect 1044 85585 1068 85641
rect 1124 85585 1148 85641
rect 1044 85517 1148 85585
rect 1044 85461 1068 85517
rect 1124 85461 1148 85517
rect 1044 85393 1148 85461
rect 1044 85337 1068 85393
rect 1124 85337 1148 85393
rect 1044 85269 1148 85337
rect 1044 85213 1068 85269
rect 1124 85213 1148 85269
rect 1044 85145 1148 85213
rect 1044 85089 1068 85145
rect 1124 85089 1148 85145
rect 1044 85021 1148 85089
rect 1044 84965 1068 85021
rect 1124 84965 1148 85021
rect 1044 84897 1148 84965
rect 1044 84841 1068 84897
rect 1124 84841 1148 84897
rect 1044 84773 1148 84841
rect 1044 84717 1068 84773
rect 1124 84717 1148 84773
rect 1044 84649 1148 84717
rect 1044 84593 1068 84649
rect 1124 84593 1148 84649
rect 1044 84525 1148 84593
rect 1044 84469 1068 84525
rect 1124 84469 1148 84525
rect 1044 84401 1148 84469
rect 1044 84345 1068 84401
rect 1124 84345 1148 84401
rect 1044 84277 1148 84345
rect 1044 84221 1068 84277
rect 1124 84221 1148 84277
rect 1044 84153 1148 84221
rect 1044 84097 1068 84153
rect 1124 84097 1148 84153
rect 1044 84029 1148 84097
rect 1044 83973 1068 84029
rect 1124 83973 1148 84029
rect 1044 83905 1148 83973
rect 1044 83849 1068 83905
rect 1124 83849 1148 83905
rect 1044 83798 1148 83849
rect 1168 85889 1644 85940
rect 1168 85833 1192 85889
rect 1248 85833 1316 85889
rect 1372 85833 1440 85889
rect 1496 85833 1564 85889
rect 1620 85833 1644 85889
rect 1168 85765 1644 85833
rect 1168 85709 1192 85765
rect 1248 85709 1316 85765
rect 1372 85709 1440 85765
rect 1496 85709 1564 85765
rect 1620 85709 1644 85765
rect 1168 85641 1644 85709
rect 1168 85585 1192 85641
rect 1248 85585 1316 85641
rect 1372 85585 1440 85641
rect 1496 85585 1564 85641
rect 1620 85585 1644 85641
rect 1168 85517 1644 85585
rect 1168 85461 1192 85517
rect 1248 85461 1316 85517
rect 1372 85461 1440 85517
rect 1496 85461 1564 85517
rect 1620 85461 1644 85517
rect 1168 85393 1644 85461
rect 1168 85337 1192 85393
rect 1248 85337 1316 85393
rect 1372 85337 1440 85393
rect 1496 85337 1564 85393
rect 1620 85337 1644 85393
rect 1168 85269 1644 85337
rect 1168 85213 1192 85269
rect 1248 85213 1316 85269
rect 1372 85213 1440 85269
rect 1496 85213 1564 85269
rect 1620 85213 1644 85269
rect 1168 85145 1644 85213
rect 1168 85089 1192 85145
rect 1248 85089 1316 85145
rect 1372 85089 1440 85145
rect 1496 85089 1564 85145
rect 1620 85089 1644 85145
rect 1168 85021 1644 85089
rect 1168 84965 1192 85021
rect 1248 84965 1316 85021
rect 1372 84965 1440 85021
rect 1496 84965 1564 85021
rect 1620 84965 1644 85021
rect 1168 84897 1644 84965
rect 1168 84841 1192 84897
rect 1248 84841 1316 84897
rect 1372 84841 1440 84897
rect 1496 84841 1564 84897
rect 1620 84841 1644 84897
rect 1168 84773 1644 84841
rect 1168 84717 1192 84773
rect 1248 84717 1316 84773
rect 1372 84717 1440 84773
rect 1496 84717 1564 84773
rect 1620 84717 1644 84773
rect 1168 84649 1644 84717
rect 1168 84593 1192 84649
rect 1248 84593 1316 84649
rect 1372 84593 1440 84649
rect 1496 84593 1564 84649
rect 1620 84593 1644 84649
rect 1168 84525 1644 84593
rect 1168 84469 1192 84525
rect 1248 84469 1316 84525
rect 1372 84469 1440 84525
rect 1496 84469 1564 84525
rect 1620 84469 1644 84525
rect 1168 84401 1644 84469
rect 1168 84345 1192 84401
rect 1248 84345 1316 84401
rect 1372 84345 1440 84401
rect 1496 84345 1564 84401
rect 1620 84345 1644 84401
rect 1168 84277 1644 84345
rect 1168 84221 1192 84277
rect 1248 84221 1316 84277
rect 1372 84221 1440 84277
rect 1496 84221 1564 84277
rect 1620 84221 1644 84277
rect 1168 84153 1644 84221
rect 1168 84097 1192 84153
rect 1248 84097 1316 84153
rect 1372 84097 1440 84153
rect 1496 84097 1564 84153
rect 1620 84097 1644 84153
rect 1168 84029 1644 84097
rect 1168 83973 1192 84029
rect 1248 83973 1316 84029
rect 1372 83973 1440 84029
rect 1496 83973 1564 84029
rect 1620 83973 1644 84029
rect 1168 83905 1644 83973
rect 1168 83849 1192 83905
rect 1248 83849 1316 83905
rect 1372 83849 1440 83905
rect 1496 83849 1564 83905
rect 1620 83849 1644 83905
rect 1168 83798 1644 83849
rect 85726 85889 85830 85940
rect 85726 85833 85750 85889
rect 85806 85833 85830 85889
rect 85726 85765 85830 85833
rect 85726 85709 85750 85765
rect 85806 85709 85830 85765
rect 85726 85641 85830 85709
rect 85726 85585 85750 85641
rect 85806 85585 85830 85641
rect 85726 85517 85830 85585
rect 85726 85461 85750 85517
rect 85806 85461 85830 85517
rect 85726 85393 85830 85461
rect 85726 85337 85750 85393
rect 85806 85337 85830 85393
rect 85726 85269 85830 85337
rect 85726 85213 85750 85269
rect 85806 85213 85830 85269
rect 85726 85145 85830 85213
rect 85726 85089 85750 85145
rect 85806 85089 85830 85145
rect 85726 85021 85830 85089
rect 85726 84965 85750 85021
rect 85806 84965 85830 85021
rect 85726 84897 85830 84965
rect 85726 84841 85750 84897
rect 85806 84841 85830 84897
rect 85726 84773 85830 84841
rect 85726 84717 85750 84773
rect 85806 84717 85830 84773
rect 85726 84649 85830 84717
rect 85726 84593 85750 84649
rect 85806 84593 85830 84649
rect 85726 84525 85830 84593
rect 85726 84469 85750 84525
rect 85806 84469 85830 84525
rect 85726 84401 85830 84469
rect 85726 84345 85750 84401
rect 85806 84345 85830 84401
rect 85726 84277 85830 84345
rect 85726 84221 85750 84277
rect 85806 84221 85830 84277
rect 85726 84153 85830 84221
rect 85726 84097 85750 84153
rect 85806 84097 85830 84153
rect 85726 84029 85830 84097
rect 85726 83973 85750 84029
rect 85806 83973 85830 84029
rect 85726 83905 85830 83973
rect 85726 83849 85750 83905
rect 85806 83849 85830 83905
rect 85726 83798 85830 83849
rect 85850 85889 86326 85940
rect 85850 85833 85874 85889
rect 85930 85833 85998 85889
rect 86054 85833 86122 85889
rect 86178 85833 86246 85889
rect 86302 85833 86326 85889
rect 85850 85765 86326 85833
rect 85850 85709 85874 85765
rect 85930 85709 85998 85765
rect 86054 85709 86122 85765
rect 86178 85709 86246 85765
rect 86302 85709 86326 85765
rect 85850 85641 86326 85709
rect 85850 85585 85874 85641
rect 85930 85585 85998 85641
rect 86054 85585 86122 85641
rect 86178 85585 86246 85641
rect 86302 85585 86326 85641
rect 85850 85517 86326 85585
rect 85850 85461 85874 85517
rect 85930 85461 85998 85517
rect 86054 85461 86122 85517
rect 86178 85461 86246 85517
rect 86302 85461 86326 85517
rect 85850 85393 86326 85461
rect 85850 85337 85874 85393
rect 85930 85337 85998 85393
rect 86054 85337 86122 85393
rect 86178 85337 86246 85393
rect 86302 85337 86326 85393
rect 85850 85269 86326 85337
rect 85850 85213 85874 85269
rect 85930 85213 85998 85269
rect 86054 85213 86122 85269
rect 86178 85213 86246 85269
rect 86302 85213 86326 85269
rect 85850 85145 86326 85213
rect 85850 85089 85874 85145
rect 85930 85089 85998 85145
rect 86054 85089 86122 85145
rect 86178 85089 86246 85145
rect 86302 85089 86326 85145
rect 85850 85021 86326 85089
rect 85850 84965 85874 85021
rect 85930 84965 85998 85021
rect 86054 84965 86122 85021
rect 86178 84965 86246 85021
rect 86302 84965 86326 85021
rect 85850 84897 86326 84965
rect 85850 84841 85874 84897
rect 85930 84841 85998 84897
rect 86054 84841 86122 84897
rect 86178 84841 86246 84897
rect 86302 84841 86326 84897
rect 85850 84773 86326 84841
rect 85850 84717 85874 84773
rect 85930 84717 85998 84773
rect 86054 84717 86122 84773
rect 86178 84717 86246 84773
rect 86302 84717 86326 84773
rect 85850 84649 86326 84717
rect 85850 84593 85874 84649
rect 85930 84593 85998 84649
rect 86054 84593 86122 84649
rect 86178 84593 86246 84649
rect 86302 84593 86326 84649
rect 85850 84525 86326 84593
rect 85850 84469 85874 84525
rect 85930 84469 85998 84525
rect 86054 84469 86122 84525
rect 86178 84469 86246 84525
rect 86302 84469 86326 84525
rect 85850 84401 86326 84469
rect 85850 84345 85874 84401
rect 85930 84345 85998 84401
rect 86054 84345 86122 84401
rect 86178 84345 86246 84401
rect 86302 84345 86326 84401
rect 85850 84277 86326 84345
rect 85850 84221 85874 84277
rect 85930 84221 85998 84277
rect 86054 84221 86122 84277
rect 86178 84221 86246 84277
rect 86302 84221 86326 84277
rect 85850 84153 86326 84221
rect 85850 84097 85874 84153
rect 85930 84097 85998 84153
rect 86054 84097 86122 84153
rect 86178 84097 86246 84153
rect 86302 84097 86326 84153
rect 85850 84029 86326 84097
rect 85850 83973 85874 84029
rect 85930 83973 85998 84029
rect 86054 83973 86122 84029
rect 86178 83973 86246 84029
rect 86302 83973 86326 84029
rect 85850 83905 86326 83973
rect 85850 83849 85874 83905
rect 85930 83849 85998 83905
rect 86054 83849 86122 83905
rect 86178 83849 86246 83905
rect 86302 83849 86326 83905
rect 85850 83798 86326 83849
rect 1844 83587 1948 83648
rect 1844 83531 1868 83587
rect 1924 83531 1948 83587
rect 1844 83463 1948 83531
rect 1844 83407 1868 83463
rect 1924 83407 1948 83463
rect 1844 83339 1948 83407
rect 1844 83283 1868 83339
rect 1924 83283 1948 83339
rect 1844 83215 1948 83283
rect 1844 83159 1868 83215
rect 1924 83159 1948 83215
rect 1844 83091 1948 83159
rect 1844 83035 1868 83091
rect 1924 83035 1948 83091
rect 1844 82967 1948 83035
rect 1844 82911 1868 82967
rect 1924 82911 1948 82967
rect 1844 82843 1948 82911
rect 1844 82787 1868 82843
rect 1924 82787 1948 82843
rect 1844 82719 1948 82787
rect 1844 82663 1868 82719
rect 1924 82663 1948 82719
rect 1844 82595 1948 82663
rect 1844 82539 1868 82595
rect 1924 82539 1948 82595
rect 1844 82471 1948 82539
rect 1844 82415 1868 82471
rect 1924 82415 1948 82471
rect 1844 82347 1948 82415
rect 1844 82291 1868 82347
rect 1924 82291 1948 82347
rect 1844 82223 1948 82291
rect 1844 82167 1868 82223
rect 1924 82167 1948 82223
rect 1844 82099 1948 82167
rect 1844 82043 1868 82099
rect 1924 82043 1948 82099
rect 1844 81975 1948 82043
rect 1844 81919 1868 81975
rect 1924 81919 1948 81975
rect 1844 81851 1948 81919
rect 1844 81795 1868 81851
rect 1924 81795 1948 81851
rect 1844 81727 1948 81795
rect 1844 81671 1868 81727
rect 1924 81671 1948 81727
rect 1844 81603 1948 81671
rect 1844 81547 1868 81603
rect 1924 81547 1948 81603
rect 1844 81479 1948 81547
rect 1844 81423 1868 81479
rect 1924 81423 1948 81479
rect 1844 81355 1948 81423
rect 1844 81299 1868 81355
rect 1924 81299 1948 81355
rect 1844 81231 1948 81299
rect 1844 81175 1868 81231
rect 1924 81175 1948 81231
rect 1844 81107 1948 81175
rect 1844 81051 1868 81107
rect 1924 81051 1948 81107
rect 1844 80983 1948 81051
rect 1844 80927 1868 80983
rect 1924 80927 1948 80983
rect 1844 80859 1948 80927
rect 1844 80803 1868 80859
rect 1924 80803 1948 80859
rect 1844 80735 1948 80803
rect 1844 80679 1868 80735
rect 1924 80679 1948 80735
rect 1844 80611 1948 80679
rect 1844 80555 1868 80611
rect 1924 80555 1948 80611
rect 1844 80487 1948 80555
rect 1844 80431 1868 80487
rect 1924 80431 1948 80487
rect 1844 80363 1948 80431
rect 1844 80307 1868 80363
rect 1924 80307 1948 80363
rect 1844 80246 1948 80307
rect 1968 83587 2444 83648
rect 1968 83531 1992 83587
rect 2048 83531 2116 83587
rect 2172 83531 2240 83587
rect 2296 83531 2364 83587
rect 2420 83531 2444 83587
rect 1968 83463 2444 83531
rect 1968 83407 1992 83463
rect 2048 83407 2116 83463
rect 2172 83407 2240 83463
rect 2296 83407 2364 83463
rect 2420 83407 2444 83463
rect 1968 83339 2444 83407
rect 1968 83283 1992 83339
rect 2048 83283 2116 83339
rect 2172 83283 2240 83339
rect 2296 83283 2364 83339
rect 2420 83283 2444 83339
rect 1968 83215 2444 83283
rect 1968 83159 1992 83215
rect 2048 83159 2116 83215
rect 2172 83159 2240 83215
rect 2296 83159 2364 83215
rect 2420 83159 2444 83215
rect 1968 83091 2444 83159
rect 1968 83035 1992 83091
rect 2048 83035 2116 83091
rect 2172 83035 2240 83091
rect 2296 83035 2364 83091
rect 2420 83035 2444 83091
rect 1968 82967 2444 83035
rect 1968 82911 1992 82967
rect 2048 82911 2116 82967
rect 2172 82911 2240 82967
rect 2296 82911 2364 82967
rect 2420 82911 2444 82967
rect 1968 82843 2444 82911
rect 1968 82787 1992 82843
rect 2048 82787 2116 82843
rect 2172 82787 2240 82843
rect 2296 82787 2364 82843
rect 2420 82787 2444 82843
rect 1968 82719 2444 82787
rect 1968 82663 1992 82719
rect 2048 82663 2116 82719
rect 2172 82663 2240 82719
rect 2296 82663 2364 82719
rect 2420 82663 2444 82719
rect 1968 82595 2444 82663
rect 1968 82539 1992 82595
rect 2048 82539 2116 82595
rect 2172 82539 2240 82595
rect 2296 82539 2364 82595
rect 2420 82539 2444 82595
rect 1968 82471 2444 82539
rect 1968 82415 1992 82471
rect 2048 82415 2116 82471
rect 2172 82415 2240 82471
rect 2296 82415 2364 82471
rect 2420 82415 2444 82471
rect 1968 82347 2444 82415
rect 1968 82291 1992 82347
rect 2048 82291 2116 82347
rect 2172 82291 2240 82347
rect 2296 82291 2364 82347
rect 2420 82291 2444 82347
rect 1968 82223 2444 82291
rect 1968 82167 1992 82223
rect 2048 82167 2116 82223
rect 2172 82167 2240 82223
rect 2296 82167 2364 82223
rect 2420 82167 2444 82223
rect 1968 82099 2444 82167
rect 1968 82043 1992 82099
rect 2048 82043 2116 82099
rect 2172 82043 2240 82099
rect 2296 82043 2364 82099
rect 2420 82043 2444 82099
rect 1968 81975 2444 82043
rect 1968 81919 1992 81975
rect 2048 81919 2116 81975
rect 2172 81919 2240 81975
rect 2296 81919 2364 81975
rect 2420 81919 2444 81975
rect 1968 81851 2444 81919
rect 1968 81795 1992 81851
rect 2048 81795 2116 81851
rect 2172 81795 2240 81851
rect 2296 81795 2364 81851
rect 2420 81795 2444 81851
rect 1968 81727 2444 81795
rect 1968 81671 1992 81727
rect 2048 81671 2116 81727
rect 2172 81671 2240 81727
rect 2296 81671 2364 81727
rect 2420 81671 2444 81727
rect 1968 81603 2444 81671
rect 1968 81547 1992 81603
rect 2048 81547 2116 81603
rect 2172 81547 2240 81603
rect 2296 81547 2364 81603
rect 2420 81547 2444 81603
rect 1968 81479 2444 81547
rect 1968 81423 1992 81479
rect 2048 81423 2116 81479
rect 2172 81423 2240 81479
rect 2296 81423 2364 81479
rect 2420 81423 2444 81479
rect 1968 81355 2444 81423
rect 1968 81299 1992 81355
rect 2048 81299 2116 81355
rect 2172 81299 2240 81355
rect 2296 81299 2364 81355
rect 2420 81299 2444 81355
rect 1968 81231 2444 81299
rect 1968 81175 1992 81231
rect 2048 81175 2116 81231
rect 2172 81175 2240 81231
rect 2296 81175 2364 81231
rect 2420 81175 2444 81231
rect 1968 81107 2444 81175
rect 1968 81051 1992 81107
rect 2048 81051 2116 81107
rect 2172 81051 2240 81107
rect 2296 81051 2364 81107
rect 2420 81051 2444 81107
rect 1968 80983 2444 81051
rect 1968 80927 1992 80983
rect 2048 80927 2116 80983
rect 2172 80927 2240 80983
rect 2296 80927 2364 80983
rect 2420 80927 2444 80983
rect 1968 80859 2444 80927
rect 1968 80803 1992 80859
rect 2048 80803 2116 80859
rect 2172 80803 2240 80859
rect 2296 80803 2364 80859
rect 2420 80803 2444 80859
rect 1968 80735 2444 80803
rect 1968 80679 1992 80735
rect 2048 80679 2116 80735
rect 2172 80679 2240 80735
rect 2296 80679 2364 80735
rect 2420 80679 2444 80735
rect 1968 80611 2444 80679
rect 1968 80555 1992 80611
rect 2048 80555 2116 80611
rect 2172 80555 2240 80611
rect 2296 80555 2364 80611
rect 2420 80555 2444 80611
rect 1968 80487 2444 80555
rect 1968 80431 1992 80487
rect 2048 80431 2116 80487
rect 2172 80431 2240 80487
rect 2296 80431 2364 80487
rect 2420 80431 2444 80487
rect 1968 80363 2444 80431
rect 1968 80307 1992 80363
rect 2048 80307 2116 80363
rect 2172 80307 2240 80363
rect 2296 80307 2364 80363
rect 2420 80307 2444 80363
rect 1968 80246 2444 80307
rect 86526 83587 86630 83648
rect 86526 83531 86550 83587
rect 86606 83531 86630 83587
rect 86526 83463 86630 83531
rect 86526 83407 86550 83463
rect 86606 83407 86630 83463
rect 86526 83339 86630 83407
rect 86526 83283 86550 83339
rect 86606 83283 86630 83339
rect 86526 83215 86630 83283
rect 86526 83159 86550 83215
rect 86606 83159 86630 83215
rect 86526 83091 86630 83159
rect 86526 83035 86550 83091
rect 86606 83035 86630 83091
rect 86526 82967 86630 83035
rect 86526 82911 86550 82967
rect 86606 82911 86630 82967
rect 86526 82843 86630 82911
rect 86526 82787 86550 82843
rect 86606 82787 86630 82843
rect 86526 82719 86630 82787
rect 86526 82663 86550 82719
rect 86606 82663 86630 82719
rect 86526 82595 86630 82663
rect 86526 82539 86550 82595
rect 86606 82539 86630 82595
rect 86526 82471 86630 82539
rect 86526 82415 86550 82471
rect 86606 82415 86630 82471
rect 86526 82347 86630 82415
rect 86526 82291 86550 82347
rect 86606 82291 86630 82347
rect 86526 82223 86630 82291
rect 86526 82167 86550 82223
rect 86606 82167 86630 82223
rect 86526 82099 86630 82167
rect 86526 82043 86550 82099
rect 86606 82043 86630 82099
rect 86526 81975 86630 82043
rect 86526 81919 86550 81975
rect 86606 81919 86630 81975
rect 86526 81851 86630 81919
rect 86526 81795 86550 81851
rect 86606 81795 86630 81851
rect 86526 81727 86630 81795
rect 86526 81671 86550 81727
rect 86606 81671 86630 81727
rect 86526 81603 86630 81671
rect 86526 81547 86550 81603
rect 86606 81547 86630 81603
rect 86526 81479 86630 81547
rect 86526 81423 86550 81479
rect 86606 81423 86630 81479
rect 86526 81355 86630 81423
rect 86526 81299 86550 81355
rect 86606 81299 86630 81355
rect 86526 81231 86630 81299
rect 86526 81175 86550 81231
rect 86606 81175 86630 81231
rect 86526 81107 86630 81175
rect 86526 81051 86550 81107
rect 86606 81051 86630 81107
rect 86526 80983 86630 81051
rect 86526 80927 86550 80983
rect 86606 80927 86630 80983
rect 86526 80859 86630 80927
rect 86526 80803 86550 80859
rect 86606 80803 86630 80859
rect 86526 80735 86630 80803
rect 86526 80679 86550 80735
rect 86606 80679 86630 80735
rect 86526 80611 86630 80679
rect 86526 80555 86550 80611
rect 86606 80555 86630 80611
rect 86526 80487 86630 80555
rect 86526 80431 86550 80487
rect 86606 80431 86630 80487
rect 86526 80363 86630 80431
rect 86526 80307 86550 80363
rect 86606 80307 86630 80363
rect 86526 80246 86630 80307
rect 86650 83587 87126 83648
rect 86650 83531 86674 83587
rect 86730 83531 86798 83587
rect 86854 83531 86922 83587
rect 86978 83531 87046 83587
rect 87102 83531 87126 83587
rect 86650 83463 87126 83531
rect 86650 83407 86674 83463
rect 86730 83407 86798 83463
rect 86854 83407 86922 83463
rect 86978 83407 87046 83463
rect 87102 83407 87126 83463
rect 86650 83339 87126 83407
rect 86650 83283 86674 83339
rect 86730 83283 86798 83339
rect 86854 83283 86922 83339
rect 86978 83283 87046 83339
rect 87102 83283 87126 83339
rect 86650 83215 87126 83283
rect 86650 83159 86674 83215
rect 86730 83159 86798 83215
rect 86854 83159 86922 83215
rect 86978 83159 87046 83215
rect 87102 83159 87126 83215
rect 86650 83091 87126 83159
rect 86650 83035 86674 83091
rect 86730 83035 86798 83091
rect 86854 83035 86922 83091
rect 86978 83035 87046 83091
rect 87102 83035 87126 83091
rect 86650 82967 87126 83035
rect 86650 82911 86674 82967
rect 86730 82911 86798 82967
rect 86854 82911 86922 82967
rect 86978 82911 87046 82967
rect 87102 82911 87126 82967
rect 86650 82843 87126 82911
rect 86650 82787 86674 82843
rect 86730 82787 86798 82843
rect 86854 82787 86922 82843
rect 86978 82787 87046 82843
rect 87102 82787 87126 82843
rect 86650 82719 87126 82787
rect 86650 82663 86674 82719
rect 86730 82663 86798 82719
rect 86854 82663 86922 82719
rect 86978 82663 87046 82719
rect 87102 82663 87126 82719
rect 86650 82595 87126 82663
rect 86650 82539 86674 82595
rect 86730 82539 86798 82595
rect 86854 82539 86922 82595
rect 86978 82539 87046 82595
rect 87102 82539 87126 82595
rect 86650 82471 87126 82539
rect 86650 82415 86674 82471
rect 86730 82415 86798 82471
rect 86854 82415 86922 82471
rect 86978 82415 87046 82471
rect 87102 82415 87126 82471
rect 86650 82347 87126 82415
rect 86650 82291 86674 82347
rect 86730 82291 86798 82347
rect 86854 82291 86922 82347
rect 86978 82291 87046 82347
rect 87102 82291 87126 82347
rect 86650 82223 87126 82291
rect 86650 82167 86674 82223
rect 86730 82167 86798 82223
rect 86854 82167 86922 82223
rect 86978 82167 87046 82223
rect 87102 82167 87126 82223
rect 86650 82099 87126 82167
rect 86650 82043 86674 82099
rect 86730 82043 86798 82099
rect 86854 82043 86922 82099
rect 86978 82043 87046 82099
rect 87102 82043 87126 82099
rect 86650 81975 87126 82043
rect 86650 81919 86674 81975
rect 86730 81919 86798 81975
rect 86854 81919 86922 81975
rect 86978 81919 87046 81975
rect 87102 81919 87126 81975
rect 86650 81851 87126 81919
rect 86650 81795 86674 81851
rect 86730 81795 86798 81851
rect 86854 81795 86922 81851
rect 86978 81795 87046 81851
rect 87102 81795 87126 81851
rect 86650 81727 87126 81795
rect 86650 81671 86674 81727
rect 86730 81671 86798 81727
rect 86854 81671 86922 81727
rect 86978 81671 87046 81727
rect 87102 81671 87126 81727
rect 86650 81603 87126 81671
rect 86650 81547 86674 81603
rect 86730 81547 86798 81603
rect 86854 81547 86922 81603
rect 86978 81547 87046 81603
rect 87102 81547 87126 81603
rect 86650 81479 87126 81547
rect 86650 81423 86674 81479
rect 86730 81423 86798 81479
rect 86854 81423 86922 81479
rect 86978 81423 87046 81479
rect 87102 81423 87126 81479
rect 86650 81355 87126 81423
rect 86650 81299 86674 81355
rect 86730 81299 86798 81355
rect 86854 81299 86922 81355
rect 86978 81299 87046 81355
rect 87102 81299 87126 81355
rect 86650 81231 87126 81299
rect 86650 81175 86674 81231
rect 86730 81175 86798 81231
rect 86854 81175 86922 81231
rect 86978 81175 87046 81231
rect 87102 81175 87126 81231
rect 86650 81107 87126 81175
rect 86650 81051 86674 81107
rect 86730 81051 86798 81107
rect 86854 81051 86922 81107
rect 86978 81051 87046 81107
rect 87102 81051 87126 81107
rect 86650 80983 87126 81051
rect 86650 80927 86674 80983
rect 86730 80927 86798 80983
rect 86854 80927 86922 80983
rect 86978 80927 87046 80983
rect 87102 80927 87126 80983
rect 86650 80859 87126 80927
rect 86650 80803 86674 80859
rect 86730 80803 86798 80859
rect 86854 80803 86922 80859
rect 86978 80803 87046 80859
rect 87102 80803 87126 80859
rect 86650 80735 87126 80803
rect 86650 80679 86674 80735
rect 86730 80679 86798 80735
rect 86854 80679 86922 80735
rect 86978 80679 87046 80735
rect 87102 80679 87126 80735
rect 86650 80611 87126 80679
rect 86650 80555 86674 80611
rect 86730 80555 86798 80611
rect 86854 80555 86922 80611
rect 86978 80555 87046 80611
rect 87102 80555 87126 80611
rect 86650 80487 87126 80555
rect 86650 80431 86674 80487
rect 86730 80431 86798 80487
rect 86854 80431 86922 80487
rect 86978 80431 87046 80487
rect 87102 80431 87126 80487
rect 86650 80363 87126 80431
rect 86650 80307 86674 80363
rect 86730 80307 86798 80363
rect 86854 80307 86922 80363
rect 86978 80307 87046 80363
rect 87102 80307 87126 80363
rect 86650 80246 87126 80307
rect 86526 76656 86630 76694
rect 86526 76600 86550 76656
rect 86606 76600 86630 76656
rect 86526 76532 86630 76600
rect 86526 76476 86550 76532
rect 86606 76476 86630 76532
rect 86526 76408 86630 76476
rect 86526 76352 86550 76408
rect 86606 76352 86630 76408
rect 86526 76284 86630 76352
rect 86526 76228 86550 76284
rect 86606 76228 86630 76284
rect 86526 76160 86630 76228
rect 86526 76104 86550 76160
rect 86606 76104 86630 76160
rect 86526 76036 86630 76104
rect 86526 75980 86550 76036
rect 86606 75980 86630 76036
rect 86526 75912 86630 75980
rect 86526 75856 86550 75912
rect 86606 75856 86630 75912
rect 86526 75788 86630 75856
rect 86526 75732 86550 75788
rect 86606 75732 86630 75788
rect 86526 75694 86630 75732
rect 86650 76656 87126 76694
rect 86650 76600 86674 76656
rect 86730 76600 86798 76656
rect 86854 76600 86922 76656
rect 86978 76600 87046 76656
rect 87102 76600 87126 76656
rect 86650 76532 87126 76600
rect 86650 76476 86674 76532
rect 86730 76476 86798 76532
rect 86854 76476 86922 76532
rect 86978 76476 87046 76532
rect 87102 76476 87126 76532
rect 86650 76408 87126 76476
rect 86650 76352 86674 76408
rect 86730 76352 86798 76408
rect 86854 76352 86922 76408
rect 86978 76352 87046 76408
rect 87102 76352 87126 76408
rect 86650 76284 87126 76352
rect 86650 76228 86674 76284
rect 86730 76228 86798 76284
rect 86854 76228 86922 76284
rect 86978 76228 87046 76284
rect 87102 76228 87126 76284
rect 86650 76160 87126 76228
rect 86650 76104 86674 76160
rect 86730 76104 86798 76160
rect 86854 76104 86922 76160
rect 86978 76104 87046 76160
rect 87102 76104 87126 76160
rect 86650 76036 87126 76104
rect 86650 75980 86674 76036
rect 86730 75980 86798 76036
rect 86854 75980 86922 76036
rect 86978 75980 87046 76036
rect 87102 75980 87126 76036
rect 86650 75912 87126 75980
rect 86650 75856 86674 75912
rect 86730 75856 86798 75912
rect 86854 75856 86922 75912
rect 86978 75856 87046 75912
rect 87102 75856 87126 75912
rect 86650 75788 87126 75856
rect 86650 75732 86674 75788
rect 86730 75732 86798 75788
rect 86854 75732 86922 75788
rect 86978 75732 87046 75788
rect 87102 75732 87126 75788
rect 86650 75694 87126 75732
rect 1044 75000 1148 75038
rect 1044 74944 1068 75000
rect 1124 74944 1148 75000
rect 1044 74876 1148 74944
rect 1044 74820 1068 74876
rect 1124 74820 1148 74876
rect 1044 74752 1148 74820
rect 1044 74696 1068 74752
rect 1124 74696 1148 74752
rect 1044 74628 1148 74696
rect 1044 74572 1068 74628
rect 1124 74572 1148 74628
rect 1044 74504 1148 74572
rect 1044 74448 1068 74504
rect 1124 74448 1148 74504
rect 1044 74380 1148 74448
rect 1044 74324 1068 74380
rect 1124 74324 1148 74380
rect 1044 74256 1148 74324
rect 1044 74200 1068 74256
rect 1124 74200 1148 74256
rect 1044 74132 1148 74200
rect 1044 74076 1068 74132
rect 1124 74076 1148 74132
rect 1044 74038 1148 74076
rect 1168 75000 1644 75038
rect 1168 74944 1192 75000
rect 1248 74944 1316 75000
rect 1372 74944 1440 75000
rect 1496 74944 1564 75000
rect 1620 74944 1644 75000
rect 1168 74876 1644 74944
rect 1168 74820 1192 74876
rect 1248 74820 1316 74876
rect 1372 74820 1440 74876
rect 1496 74820 1564 74876
rect 1620 74820 1644 74876
rect 1168 74752 1644 74820
rect 1168 74696 1192 74752
rect 1248 74696 1316 74752
rect 1372 74696 1440 74752
rect 1496 74696 1564 74752
rect 1620 74696 1644 74752
rect 1168 74628 1644 74696
rect 1168 74572 1192 74628
rect 1248 74572 1316 74628
rect 1372 74572 1440 74628
rect 1496 74572 1564 74628
rect 1620 74572 1644 74628
rect 1168 74504 1644 74572
rect 1168 74448 1192 74504
rect 1248 74448 1316 74504
rect 1372 74448 1440 74504
rect 1496 74448 1564 74504
rect 1620 74448 1644 74504
rect 1168 74380 1644 74448
rect 1168 74324 1192 74380
rect 1248 74324 1316 74380
rect 1372 74324 1440 74380
rect 1496 74324 1564 74380
rect 1620 74324 1644 74380
rect 1168 74256 1644 74324
rect 1168 74200 1192 74256
rect 1248 74200 1316 74256
rect 1372 74200 1440 74256
rect 1496 74200 1564 74256
rect 1620 74200 1644 74256
rect 1168 74132 1644 74200
rect 1168 74076 1192 74132
rect 1248 74076 1316 74132
rect 1372 74076 1440 74132
rect 1496 74076 1564 74132
rect 1620 74076 1644 74132
rect 1168 74038 1644 74076
rect 85726 75000 85830 75038
rect 85726 74944 85750 75000
rect 85806 74944 85830 75000
rect 85726 74876 85830 74944
rect 85726 74820 85750 74876
rect 85806 74820 85830 74876
rect 85726 74752 85830 74820
rect 85726 74696 85750 74752
rect 85806 74696 85830 74752
rect 85726 74628 85830 74696
rect 85726 74572 85750 74628
rect 85806 74572 85830 74628
rect 85726 74504 85830 74572
rect 85726 74448 85750 74504
rect 85806 74448 85830 74504
rect 85726 74380 85830 74448
rect 85726 74324 85750 74380
rect 85806 74324 85830 74380
rect 85726 74256 85830 74324
rect 85726 74200 85750 74256
rect 85806 74200 85830 74256
rect 85726 74132 85830 74200
rect 85726 74076 85750 74132
rect 85806 74076 85830 74132
rect 85726 74038 85830 74076
rect 85850 75000 86326 75038
rect 85850 74944 85874 75000
rect 85930 74944 85998 75000
rect 86054 74944 86122 75000
rect 86178 74944 86246 75000
rect 86302 74944 86326 75000
rect 85850 74876 86326 74944
rect 85850 74820 85874 74876
rect 85930 74820 85998 74876
rect 86054 74820 86122 74876
rect 86178 74820 86246 74876
rect 86302 74820 86326 74876
rect 85850 74752 86326 74820
rect 85850 74696 85874 74752
rect 85930 74696 85998 74752
rect 86054 74696 86122 74752
rect 86178 74696 86246 74752
rect 86302 74696 86326 74752
rect 85850 74628 86326 74696
rect 85850 74572 85874 74628
rect 85930 74572 85998 74628
rect 86054 74572 86122 74628
rect 86178 74572 86246 74628
rect 86302 74572 86326 74628
rect 85850 74504 86326 74572
rect 85850 74448 85874 74504
rect 85930 74448 85998 74504
rect 86054 74448 86122 74504
rect 86178 74448 86246 74504
rect 86302 74448 86326 74504
rect 85850 74380 86326 74448
rect 85850 74324 85874 74380
rect 85930 74324 85998 74380
rect 86054 74324 86122 74380
rect 86178 74324 86246 74380
rect 86302 74324 86326 74380
rect 85850 74256 86326 74324
rect 85850 74200 85874 74256
rect 85930 74200 85998 74256
rect 86054 74200 86122 74256
rect 86178 74200 86246 74256
rect 86302 74200 86326 74256
rect 85850 74132 86326 74200
rect 85850 74076 85874 74132
rect 85930 74076 85998 74132
rect 86054 74076 86122 74132
rect 86178 74076 86246 74132
rect 86302 74076 86326 74132
rect 85850 74038 86326 74076
rect 1906 63414 2382 63440
rect 1906 63358 1930 63414
rect 1986 63358 2054 63414
rect 2110 63358 2178 63414
rect 2234 63358 2302 63414
rect 2358 63358 2382 63414
rect 1906 63290 2382 63358
rect 1906 63234 1930 63290
rect 1986 63234 2054 63290
rect 2110 63234 2178 63290
rect 2234 63234 2302 63290
rect 2358 63234 2382 63290
rect 1906 63166 2382 63234
rect 1906 63110 1930 63166
rect 1986 63110 2054 63166
rect 2110 63110 2178 63166
rect 2234 63110 2302 63166
rect 2358 63110 2382 63166
rect 1906 63042 2382 63110
rect 1906 62986 1930 63042
rect 1986 62986 2054 63042
rect 2110 62986 2178 63042
rect 2234 62986 2302 63042
rect 2358 62986 2382 63042
rect 1906 62960 2382 62986
rect 86588 63259 87064 63316
rect 86588 63203 86612 63259
rect 86668 63203 86736 63259
rect 86792 63203 86860 63259
rect 86916 63203 86984 63259
rect 87040 63203 87064 63259
rect 86588 63135 87064 63203
rect 86588 63079 86612 63135
rect 86668 63079 86736 63135
rect 86792 63079 86860 63135
rect 86916 63079 86984 63135
rect 87040 63079 87064 63135
rect 86588 63011 87064 63079
rect 86588 62955 86612 63011
rect 86668 62955 86736 63011
rect 86792 62955 86860 63011
rect 86916 62955 86984 63011
rect 87040 62955 87064 63011
rect 86588 62887 87064 62955
rect 1906 62840 2382 62850
rect 1906 62784 1930 62840
rect 1986 62784 2054 62840
rect 2110 62784 2178 62840
rect 2234 62784 2302 62840
rect 2358 62784 2382 62840
rect 1906 62716 2382 62784
rect 86588 62831 86612 62887
rect 86668 62831 86736 62887
rect 86792 62831 86860 62887
rect 86916 62831 86984 62887
rect 87040 62831 87064 62887
rect 86588 62774 87064 62831
rect 1906 62660 1930 62716
rect 1986 62660 2054 62716
rect 2110 62660 2178 62716
rect 2234 62660 2302 62716
rect 2358 62660 2382 62716
rect 1906 62650 2382 62660
rect 1106 62064 1582 62076
rect 1106 62008 1130 62064
rect 1186 62008 1254 62064
rect 1310 62008 1378 62064
rect 1434 62008 1502 62064
rect 1558 62008 1582 62064
rect 1106 61940 1582 62008
rect 1106 61884 1130 61940
rect 1186 61884 1254 61940
rect 1310 61884 1378 61940
rect 1434 61884 1502 61940
rect 1558 61884 1582 61940
rect 1106 61816 1582 61884
rect 1106 61760 1130 61816
rect 1186 61760 1254 61816
rect 1310 61760 1378 61816
rect 1434 61760 1502 61816
rect 1558 61760 1582 61816
rect 1106 61692 1582 61760
rect 1106 61636 1130 61692
rect 1186 61636 1254 61692
rect 1310 61636 1378 61692
rect 1434 61636 1502 61692
rect 1558 61636 1582 61692
rect 1106 61624 1582 61636
rect 85788 62064 86264 62076
rect 85788 62008 85812 62064
rect 85868 62008 85936 62064
rect 85992 62008 86060 62064
rect 86116 62008 86184 62064
rect 86240 62008 86264 62064
rect 85788 61940 86264 62008
rect 85788 61884 85812 61940
rect 85868 61884 85936 61940
rect 85992 61884 86060 61940
rect 86116 61884 86184 61940
rect 86240 61884 86264 61940
rect 85788 61816 86264 61884
rect 85788 61760 85812 61816
rect 85868 61760 85936 61816
rect 85992 61760 86060 61816
rect 86116 61760 86184 61816
rect 86240 61760 86264 61816
rect 85788 61692 86264 61760
rect 85788 61636 85812 61692
rect 85868 61636 85936 61692
rect 85992 61636 86060 61692
rect 86116 61636 86184 61692
rect 86240 61636 86264 61692
rect 85788 61624 86264 61636
rect 86588 61164 87064 61176
rect 86588 61108 86612 61164
rect 86668 61108 86736 61164
rect 86792 61108 86860 61164
rect 86916 61108 86984 61164
rect 87040 61108 87064 61164
rect 1906 61040 2382 61100
rect 1906 60984 1930 61040
rect 1986 60984 2054 61040
rect 2110 60984 2178 61040
rect 2234 60984 2302 61040
rect 2358 60984 2382 61040
rect 1906 60916 2382 60984
rect 1906 60860 1930 60916
rect 1986 60860 2054 60916
rect 2110 60860 2178 60916
rect 2234 60860 2302 60916
rect 2358 60860 2382 60916
rect 1906 60800 2382 60860
rect 86588 61040 87064 61108
rect 86588 60984 86612 61040
rect 86668 60984 86736 61040
rect 86792 60984 86860 61040
rect 86916 60984 86984 61040
rect 87040 60984 87064 61040
rect 86588 60916 87064 60984
rect 86588 60860 86612 60916
rect 86668 60860 86736 60916
rect 86792 60860 86860 60916
rect 86916 60860 86984 60916
rect 87040 60860 87064 60916
rect 86588 60792 87064 60860
rect 86588 60736 86612 60792
rect 86668 60736 86736 60792
rect 86792 60736 86860 60792
rect 86916 60736 86984 60792
rect 87040 60736 87064 60792
rect 86588 60724 87064 60736
rect 1106 60264 1582 60276
rect 1106 60208 1130 60264
rect 1186 60208 1254 60264
rect 1310 60208 1378 60264
rect 1434 60208 1502 60264
rect 1558 60208 1582 60264
rect 1106 60140 1582 60208
rect 1106 60084 1130 60140
rect 1186 60084 1254 60140
rect 1310 60084 1378 60140
rect 1434 60084 1502 60140
rect 1558 60084 1582 60140
rect 1106 60016 1582 60084
rect 1106 59960 1130 60016
rect 1186 59960 1254 60016
rect 1310 59960 1378 60016
rect 1434 59960 1502 60016
rect 1558 59960 1582 60016
rect 1106 59892 1582 59960
rect 1106 59836 1130 59892
rect 1186 59836 1254 59892
rect 1310 59836 1378 59892
rect 1434 59836 1502 59892
rect 1558 59836 1582 59892
rect 1106 59824 1582 59836
rect 85788 60264 86264 60276
rect 85788 60208 85812 60264
rect 85868 60208 85936 60264
rect 85992 60208 86060 60264
rect 86116 60208 86184 60264
rect 86240 60208 86264 60264
rect 85788 60140 86264 60208
rect 85788 60084 85812 60140
rect 85868 60084 85936 60140
rect 85992 60084 86060 60140
rect 86116 60084 86184 60140
rect 86240 60084 86264 60140
rect 85788 60016 86264 60084
rect 85788 59960 85812 60016
rect 85868 59960 85936 60016
rect 85992 59960 86060 60016
rect 86116 59960 86184 60016
rect 86240 59960 86264 60016
rect 85788 59892 86264 59960
rect 85788 59836 85812 59892
rect 85868 59836 85936 59892
rect 85992 59836 86060 59892
rect 86116 59836 86184 59892
rect 86240 59836 86264 59892
rect 85788 59824 86264 59836
rect 86588 59364 87064 59376
rect 86588 59308 86612 59364
rect 86668 59308 86736 59364
rect 86792 59308 86860 59364
rect 86916 59308 86984 59364
rect 87040 59308 87064 59364
rect 1906 59240 2382 59300
rect 1906 59184 1930 59240
rect 1986 59184 2054 59240
rect 2110 59184 2178 59240
rect 2234 59184 2302 59240
rect 2358 59184 2382 59240
rect 1906 59116 2382 59184
rect 1906 59060 1930 59116
rect 1986 59060 2054 59116
rect 2110 59060 2178 59116
rect 2234 59060 2302 59116
rect 2358 59060 2382 59116
rect 1906 59000 2382 59060
rect 86588 59240 87064 59308
rect 86588 59184 86612 59240
rect 86668 59184 86736 59240
rect 86792 59184 86860 59240
rect 86916 59184 86984 59240
rect 87040 59184 87064 59240
rect 86588 59116 87064 59184
rect 86588 59060 86612 59116
rect 86668 59060 86736 59116
rect 86792 59060 86860 59116
rect 86916 59060 86984 59116
rect 87040 59060 87064 59116
rect 86588 58992 87064 59060
rect 86588 58936 86612 58992
rect 86668 58936 86736 58992
rect 86792 58936 86860 58992
rect 86916 58936 86984 58992
rect 87040 58936 87064 58992
rect 86588 58924 87064 58936
rect 1106 58464 1582 58476
rect 1106 58408 1130 58464
rect 1186 58408 1254 58464
rect 1310 58408 1378 58464
rect 1434 58408 1502 58464
rect 1558 58408 1582 58464
rect 1106 58340 1582 58408
rect 1106 58284 1130 58340
rect 1186 58284 1254 58340
rect 1310 58284 1378 58340
rect 1434 58284 1502 58340
rect 1558 58284 1582 58340
rect 1106 58216 1582 58284
rect 1106 58160 1130 58216
rect 1186 58160 1254 58216
rect 1310 58160 1378 58216
rect 1434 58160 1502 58216
rect 1558 58160 1582 58216
rect 1106 58092 1582 58160
rect 1106 58036 1130 58092
rect 1186 58036 1254 58092
rect 1310 58036 1378 58092
rect 1434 58036 1502 58092
rect 1558 58036 1582 58092
rect 1106 58024 1582 58036
rect 85788 58464 86264 58476
rect 85788 58408 85812 58464
rect 85868 58408 85936 58464
rect 85992 58408 86060 58464
rect 86116 58408 86184 58464
rect 86240 58408 86264 58464
rect 85788 58340 86264 58408
rect 85788 58284 85812 58340
rect 85868 58284 85936 58340
rect 85992 58284 86060 58340
rect 86116 58284 86184 58340
rect 86240 58284 86264 58340
rect 85788 58216 86264 58284
rect 85788 58160 85812 58216
rect 85868 58160 85936 58216
rect 85992 58160 86060 58216
rect 86116 58160 86184 58216
rect 86240 58160 86264 58216
rect 85788 58092 86264 58160
rect 85788 58036 85812 58092
rect 85868 58036 85936 58092
rect 85992 58036 86060 58092
rect 86116 58036 86184 58092
rect 86240 58036 86264 58092
rect 85788 58024 86264 58036
rect 86588 57564 87064 57576
rect 86588 57508 86612 57564
rect 86668 57508 86736 57564
rect 86792 57508 86860 57564
rect 86916 57508 86984 57564
rect 87040 57508 87064 57564
rect 1906 57440 2382 57500
rect 1906 57384 1930 57440
rect 1986 57384 2054 57440
rect 2110 57384 2178 57440
rect 2234 57384 2302 57440
rect 2358 57384 2382 57440
rect 1906 57316 2382 57384
rect 1906 57260 1930 57316
rect 1986 57260 2054 57316
rect 2110 57260 2178 57316
rect 2234 57260 2302 57316
rect 2358 57260 2382 57316
rect 1906 57200 2382 57260
rect 86588 57440 87064 57508
rect 86588 57384 86612 57440
rect 86668 57384 86736 57440
rect 86792 57384 86860 57440
rect 86916 57384 86984 57440
rect 87040 57384 87064 57440
rect 86588 57316 87064 57384
rect 86588 57260 86612 57316
rect 86668 57260 86736 57316
rect 86792 57260 86860 57316
rect 86916 57260 86984 57316
rect 87040 57260 87064 57316
rect 86588 57192 87064 57260
rect 86588 57136 86612 57192
rect 86668 57136 86736 57192
rect 86792 57136 86860 57192
rect 86916 57136 86984 57192
rect 87040 57136 87064 57192
rect 86588 57124 87064 57136
rect 1106 56664 1582 56676
rect 1106 56608 1130 56664
rect 1186 56608 1254 56664
rect 1310 56608 1378 56664
rect 1434 56608 1502 56664
rect 1558 56608 1582 56664
rect 1106 56540 1582 56608
rect 1106 56484 1130 56540
rect 1186 56484 1254 56540
rect 1310 56484 1378 56540
rect 1434 56484 1502 56540
rect 1558 56484 1582 56540
rect 1106 56416 1582 56484
rect 1106 56360 1130 56416
rect 1186 56360 1254 56416
rect 1310 56360 1378 56416
rect 1434 56360 1502 56416
rect 1558 56360 1582 56416
rect 1106 56292 1582 56360
rect 1106 56236 1130 56292
rect 1186 56236 1254 56292
rect 1310 56236 1378 56292
rect 1434 56236 1502 56292
rect 1558 56236 1582 56292
rect 1106 56224 1582 56236
rect 85788 56664 86264 56676
rect 85788 56608 85812 56664
rect 85868 56608 85936 56664
rect 85992 56608 86060 56664
rect 86116 56608 86184 56664
rect 86240 56608 86264 56664
rect 85788 56540 86264 56608
rect 85788 56484 85812 56540
rect 85868 56484 85936 56540
rect 85992 56484 86060 56540
rect 86116 56484 86184 56540
rect 86240 56484 86264 56540
rect 85788 56416 86264 56484
rect 85788 56360 85812 56416
rect 85868 56360 85936 56416
rect 85992 56360 86060 56416
rect 86116 56360 86184 56416
rect 86240 56360 86264 56416
rect 85788 56292 86264 56360
rect 85788 56236 85812 56292
rect 85868 56236 85936 56292
rect 85992 56236 86060 56292
rect 86116 56236 86184 56292
rect 86240 56236 86264 56292
rect 85788 56224 86264 56236
rect 86588 55764 87064 55776
rect 86588 55708 86612 55764
rect 86668 55708 86736 55764
rect 86792 55708 86860 55764
rect 86916 55708 86984 55764
rect 87040 55708 87064 55764
rect 1906 55640 2382 55700
rect 1906 55584 1930 55640
rect 1986 55584 2054 55640
rect 2110 55584 2178 55640
rect 2234 55584 2302 55640
rect 2358 55584 2382 55640
rect 1906 55516 2382 55584
rect 1906 55460 1930 55516
rect 1986 55460 2054 55516
rect 2110 55460 2178 55516
rect 2234 55460 2302 55516
rect 2358 55460 2382 55516
rect 1906 55400 2382 55460
rect 86588 55640 87064 55708
rect 86588 55584 86612 55640
rect 86668 55584 86736 55640
rect 86792 55584 86860 55640
rect 86916 55584 86984 55640
rect 87040 55584 87064 55640
rect 86588 55516 87064 55584
rect 86588 55460 86612 55516
rect 86668 55460 86736 55516
rect 86792 55460 86860 55516
rect 86916 55460 86984 55516
rect 87040 55460 87064 55516
rect 86588 55392 87064 55460
rect 86588 55336 86612 55392
rect 86668 55336 86736 55392
rect 86792 55336 86860 55392
rect 86916 55336 86984 55392
rect 87040 55336 87064 55392
rect 86588 55324 87064 55336
rect 1106 54864 1582 54876
rect 1106 54808 1130 54864
rect 1186 54808 1254 54864
rect 1310 54808 1378 54864
rect 1434 54808 1502 54864
rect 1558 54808 1582 54864
rect 1106 54740 1582 54808
rect 1106 54684 1130 54740
rect 1186 54684 1254 54740
rect 1310 54684 1378 54740
rect 1434 54684 1502 54740
rect 1558 54684 1582 54740
rect 1106 54616 1582 54684
rect 1106 54560 1130 54616
rect 1186 54560 1254 54616
rect 1310 54560 1378 54616
rect 1434 54560 1502 54616
rect 1558 54560 1582 54616
rect 1106 54492 1582 54560
rect 1106 54436 1130 54492
rect 1186 54436 1254 54492
rect 1310 54436 1378 54492
rect 1434 54436 1502 54492
rect 1558 54436 1582 54492
rect 1106 54424 1582 54436
rect 85788 54864 86264 54876
rect 85788 54808 85812 54864
rect 85868 54808 85936 54864
rect 85992 54808 86060 54864
rect 86116 54808 86184 54864
rect 86240 54808 86264 54864
rect 85788 54740 86264 54808
rect 85788 54684 85812 54740
rect 85868 54684 85936 54740
rect 85992 54684 86060 54740
rect 86116 54684 86184 54740
rect 86240 54684 86264 54740
rect 85788 54616 86264 54684
rect 85788 54560 85812 54616
rect 85868 54560 85936 54616
rect 85992 54560 86060 54616
rect 86116 54560 86184 54616
rect 86240 54560 86264 54616
rect 85788 54492 86264 54560
rect 85788 54436 85812 54492
rect 85868 54436 85936 54492
rect 85992 54436 86060 54492
rect 86116 54436 86184 54492
rect 86240 54436 86264 54492
rect 85788 54424 86264 54436
rect 86588 53964 87064 53976
rect 86588 53908 86612 53964
rect 86668 53908 86736 53964
rect 86792 53908 86860 53964
rect 86916 53908 86984 53964
rect 87040 53908 87064 53964
rect 1906 53840 2382 53900
rect 1906 53784 1930 53840
rect 1986 53784 2054 53840
rect 2110 53784 2178 53840
rect 2234 53784 2302 53840
rect 2358 53784 2382 53840
rect 1906 53716 2382 53784
rect 1906 53660 1930 53716
rect 1986 53660 2054 53716
rect 2110 53660 2178 53716
rect 2234 53660 2302 53716
rect 2358 53660 2382 53716
rect 1906 53600 2382 53660
rect 86588 53840 87064 53908
rect 86588 53784 86612 53840
rect 86668 53784 86736 53840
rect 86792 53784 86860 53840
rect 86916 53784 86984 53840
rect 87040 53784 87064 53840
rect 86588 53716 87064 53784
rect 86588 53660 86612 53716
rect 86668 53660 86736 53716
rect 86792 53660 86860 53716
rect 86916 53660 86984 53716
rect 87040 53660 87064 53716
rect 86588 53592 87064 53660
rect 86588 53536 86612 53592
rect 86668 53536 86736 53592
rect 86792 53536 86860 53592
rect 86916 53536 86984 53592
rect 87040 53536 87064 53592
rect 86588 53524 87064 53536
rect 1106 53064 1582 53076
rect 1106 53008 1130 53064
rect 1186 53008 1254 53064
rect 1310 53008 1378 53064
rect 1434 53008 1502 53064
rect 1558 53008 1582 53064
rect 1106 52940 1582 53008
rect 1106 52884 1130 52940
rect 1186 52884 1254 52940
rect 1310 52884 1378 52940
rect 1434 52884 1502 52940
rect 1558 52884 1582 52940
rect 1106 52816 1582 52884
rect 1106 52760 1130 52816
rect 1186 52760 1254 52816
rect 1310 52760 1378 52816
rect 1434 52760 1502 52816
rect 1558 52760 1582 52816
rect 1106 52692 1582 52760
rect 1106 52636 1130 52692
rect 1186 52636 1254 52692
rect 1310 52636 1378 52692
rect 1434 52636 1502 52692
rect 1558 52636 1582 52692
rect 1106 52624 1582 52636
rect 85788 53064 86264 53076
rect 85788 53008 85812 53064
rect 85868 53008 85936 53064
rect 85992 53008 86060 53064
rect 86116 53008 86184 53064
rect 86240 53008 86264 53064
rect 85788 52940 86264 53008
rect 85788 52884 85812 52940
rect 85868 52884 85936 52940
rect 85992 52884 86060 52940
rect 86116 52884 86184 52940
rect 86240 52884 86264 52940
rect 85788 52816 86264 52884
rect 85788 52760 85812 52816
rect 85868 52760 85936 52816
rect 85992 52760 86060 52816
rect 86116 52760 86184 52816
rect 86240 52760 86264 52816
rect 85788 52692 86264 52760
rect 85788 52636 85812 52692
rect 85868 52636 85936 52692
rect 85992 52636 86060 52692
rect 86116 52636 86184 52692
rect 86240 52636 86264 52692
rect 85788 52624 86264 52636
rect 86588 52164 87064 52176
rect 86588 52108 86612 52164
rect 86668 52108 86736 52164
rect 86792 52108 86860 52164
rect 86916 52108 86984 52164
rect 87040 52108 87064 52164
rect 1906 52040 2382 52100
rect 1906 51984 1930 52040
rect 1986 51984 2054 52040
rect 2110 51984 2178 52040
rect 2234 51984 2302 52040
rect 2358 51984 2382 52040
rect 1906 51916 2382 51984
rect 1906 51860 1930 51916
rect 1986 51860 2054 51916
rect 2110 51860 2178 51916
rect 2234 51860 2302 51916
rect 2358 51860 2382 51916
rect 1906 51800 2382 51860
rect 86588 52040 87064 52108
rect 86588 51984 86612 52040
rect 86668 51984 86736 52040
rect 86792 51984 86860 52040
rect 86916 51984 86984 52040
rect 87040 51984 87064 52040
rect 86588 51916 87064 51984
rect 86588 51860 86612 51916
rect 86668 51860 86736 51916
rect 86792 51860 86860 51916
rect 86916 51860 86984 51916
rect 87040 51860 87064 51916
rect 86588 51792 87064 51860
rect 86588 51736 86612 51792
rect 86668 51736 86736 51792
rect 86792 51736 86860 51792
rect 86916 51736 86984 51792
rect 87040 51736 87064 51792
rect 86588 51724 87064 51736
rect 1106 51264 1582 51276
rect 1106 51208 1130 51264
rect 1186 51208 1254 51264
rect 1310 51208 1378 51264
rect 1434 51208 1502 51264
rect 1558 51208 1582 51264
rect 1106 51140 1582 51208
rect 1106 51084 1130 51140
rect 1186 51084 1254 51140
rect 1310 51084 1378 51140
rect 1434 51084 1502 51140
rect 1558 51084 1582 51140
rect 1106 51016 1582 51084
rect 1106 50960 1130 51016
rect 1186 50960 1254 51016
rect 1310 50960 1378 51016
rect 1434 50960 1502 51016
rect 1558 50960 1582 51016
rect 1106 50892 1582 50960
rect 1106 50836 1130 50892
rect 1186 50836 1254 50892
rect 1310 50836 1378 50892
rect 1434 50836 1502 50892
rect 1558 50836 1582 50892
rect 1106 50824 1582 50836
rect 85788 51264 86264 51276
rect 85788 51208 85812 51264
rect 85868 51208 85936 51264
rect 85992 51208 86060 51264
rect 86116 51208 86184 51264
rect 86240 51208 86264 51264
rect 85788 51140 86264 51208
rect 85788 51084 85812 51140
rect 85868 51084 85936 51140
rect 85992 51084 86060 51140
rect 86116 51084 86184 51140
rect 86240 51084 86264 51140
rect 85788 51016 86264 51084
rect 85788 50960 85812 51016
rect 85868 50960 85936 51016
rect 85992 50960 86060 51016
rect 86116 50960 86184 51016
rect 86240 50960 86264 51016
rect 85788 50892 86264 50960
rect 85788 50836 85812 50892
rect 85868 50836 85936 50892
rect 85992 50836 86060 50892
rect 86116 50836 86184 50892
rect 86240 50836 86264 50892
rect 85788 50824 86264 50836
rect 86588 50364 87064 50376
rect 86588 50308 86612 50364
rect 86668 50308 86736 50364
rect 86792 50308 86860 50364
rect 86916 50308 86984 50364
rect 87040 50308 87064 50364
rect 1906 50240 2382 50300
rect 1906 50184 1930 50240
rect 1986 50184 2054 50240
rect 2110 50184 2178 50240
rect 2234 50184 2302 50240
rect 2358 50184 2382 50240
rect 1906 50116 2382 50184
rect 1906 50060 1930 50116
rect 1986 50060 2054 50116
rect 2110 50060 2178 50116
rect 2234 50060 2302 50116
rect 2358 50060 2382 50116
rect 1906 50000 2382 50060
rect 86588 50240 87064 50308
rect 86588 50184 86612 50240
rect 86668 50184 86736 50240
rect 86792 50184 86860 50240
rect 86916 50184 86984 50240
rect 87040 50184 87064 50240
rect 86588 50116 87064 50184
rect 86588 50060 86612 50116
rect 86668 50060 86736 50116
rect 86792 50060 86860 50116
rect 86916 50060 86984 50116
rect 87040 50060 87064 50116
rect 86588 49992 87064 50060
rect 86588 49936 86612 49992
rect 86668 49936 86736 49992
rect 86792 49936 86860 49992
rect 86916 49936 86984 49992
rect 87040 49936 87064 49992
rect 86588 49924 87064 49936
rect 1106 49464 1582 49476
rect 1106 49408 1130 49464
rect 1186 49408 1254 49464
rect 1310 49408 1378 49464
rect 1434 49408 1502 49464
rect 1558 49408 1582 49464
rect 1106 49340 1582 49408
rect 1106 49284 1130 49340
rect 1186 49284 1254 49340
rect 1310 49284 1378 49340
rect 1434 49284 1502 49340
rect 1558 49284 1582 49340
rect 1106 49216 1582 49284
rect 1106 49160 1130 49216
rect 1186 49160 1254 49216
rect 1310 49160 1378 49216
rect 1434 49160 1502 49216
rect 1558 49160 1582 49216
rect 1106 49092 1582 49160
rect 1106 49036 1130 49092
rect 1186 49036 1254 49092
rect 1310 49036 1378 49092
rect 1434 49036 1502 49092
rect 1558 49036 1582 49092
rect 1106 49024 1582 49036
rect 85788 49464 86264 49476
rect 85788 49408 85812 49464
rect 85868 49408 85936 49464
rect 85992 49408 86060 49464
rect 86116 49408 86184 49464
rect 86240 49408 86264 49464
rect 85788 49340 86264 49408
rect 85788 49284 85812 49340
rect 85868 49284 85936 49340
rect 85992 49284 86060 49340
rect 86116 49284 86184 49340
rect 86240 49284 86264 49340
rect 85788 49216 86264 49284
rect 85788 49160 85812 49216
rect 85868 49160 85936 49216
rect 85992 49160 86060 49216
rect 86116 49160 86184 49216
rect 86240 49160 86264 49216
rect 85788 49092 86264 49160
rect 85788 49036 85812 49092
rect 85868 49036 85936 49092
rect 85992 49036 86060 49092
rect 86116 49036 86184 49092
rect 86240 49036 86264 49092
rect 85788 49024 86264 49036
rect 86588 48564 87064 48576
rect 86588 48508 86612 48564
rect 86668 48508 86736 48564
rect 86792 48508 86860 48564
rect 86916 48508 86984 48564
rect 87040 48508 87064 48564
rect 1906 48440 2382 48500
rect 1906 48384 1930 48440
rect 1986 48384 2054 48440
rect 2110 48384 2178 48440
rect 2234 48384 2302 48440
rect 2358 48384 2382 48440
rect 1906 48316 2382 48384
rect 1906 48260 1930 48316
rect 1986 48260 2054 48316
rect 2110 48260 2178 48316
rect 2234 48260 2302 48316
rect 2358 48260 2382 48316
rect 1906 48200 2382 48260
rect 86588 48440 87064 48508
rect 86588 48384 86612 48440
rect 86668 48384 86736 48440
rect 86792 48384 86860 48440
rect 86916 48384 86984 48440
rect 87040 48384 87064 48440
rect 86588 48316 87064 48384
rect 86588 48260 86612 48316
rect 86668 48260 86736 48316
rect 86792 48260 86860 48316
rect 86916 48260 86984 48316
rect 87040 48260 87064 48316
rect 86588 48192 87064 48260
rect 86588 48136 86612 48192
rect 86668 48136 86736 48192
rect 86792 48136 86860 48192
rect 86916 48136 86984 48192
rect 87040 48136 87064 48192
rect 86588 48124 87064 48136
rect 1106 47664 1582 47676
rect 1106 47608 1130 47664
rect 1186 47608 1254 47664
rect 1310 47608 1378 47664
rect 1434 47608 1502 47664
rect 1558 47608 1582 47664
rect 1106 47540 1582 47608
rect 1106 47484 1130 47540
rect 1186 47484 1254 47540
rect 1310 47484 1378 47540
rect 1434 47484 1502 47540
rect 1558 47484 1582 47540
rect 1106 47416 1582 47484
rect 1106 47360 1130 47416
rect 1186 47360 1254 47416
rect 1310 47360 1378 47416
rect 1434 47360 1502 47416
rect 1558 47360 1582 47416
rect 1106 47292 1582 47360
rect 1106 47236 1130 47292
rect 1186 47236 1254 47292
rect 1310 47236 1378 47292
rect 1434 47236 1502 47292
rect 1558 47236 1582 47292
rect 1106 47224 1582 47236
rect 85788 47664 86264 47676
rect 85788 47608 85812 47664
rect 85868 47608 85936 47664
rect 85992 47608 86060 47664
rect 86116 47608 86184 47664
rect 86240 47608 86264 47664
rect 85788 47540 86264 47608
rect 85788 47484 85812 47540
rect 85868 47484 85936 47540
rect 85992 47484 86060 47540
rect 86116 47484 86184 47540
rect 86240 47484 86264 47540
rect 85788 47416 86264 47484
rect 85788 47360 85812 47416
rect 85868 47360 85936 47416
rect 85992 47360 86060 47416
rect 86116 47360 86184 47416
rect 86240 47360 86264 47416
rect 85788 47292 86264 47360
rect 85788 47236 85812 47292
rect 85868 47236 85936 47292
rect 85992 47236 86060 47292
rect 86116 47236 86184 47292
rect 86240 47236 86264 47292
rect 85788 47224 86264 47236
rect 86588 46764 87064 46776
rect 86588 46708 86612 46764
rect 86668 46708 86736 46764
rect 86792 46708 86860 46764
rect 86916 46708 86984 46764
rect 87040 46708 87064 46764
rect 1906 46640 2382 46700
rect 1906 46584 1930 46640
rect 1986 46584 2054 46640
rect 2110 46584 2178 46640
rect 2234 46584 2302 46640
rect 2358 46584 2382 46640
rect 1906 46516 2382 46584
rect 1906 46460 1930 46516
rect 1986 46460 2054 46516
rect 2110 46460 2178 46516
rect 2234 46460 2302 46516
rect 2358 46460 2382 46516
rect 1906 46400 2382 46460
rect 86588 46640 87064 46708
rect 86588 46584 86612 46640
rect 86668 46584 86736 46640
rect 86792 46584 86860 46640
rect 86916 46584 86984 46640
rect 87040 46584 87064 46640
rect 86588 46516 87064 46584
rect 86588 46460 86612 46516
rect 86668 46460 86736 46516
rect 86792 46460 86860 46516
rect 86916 46460 86984 46516
rect 87040 46460 87064 46516
rect 86588 46392 87064 46460
rect 86588 46336 86612 46392
rect 86668 46336 86736 46392
rect 86792 46336 86860 46392
rect 86916 46336 86984 46392
rect 87040 46336 87064 46392
rect 86588 46324 87064 46336
rect 1106 45864 1582 45876
rect 1106 45808 1130 45864
rect 1186 45808 1254 45864
rect 1310 45808 1378 45864
rect 1434 45808 1502 45864
rect 1558 45808 1582 45864
rect 1106 45740 1582 45808
rect 1106 45684 1130 45740
rect 1186 45684 1254 45740
rect 1310 45684 1378 45740
rect 1434 45684 1502 45740
rect 1558 45684 1582 45740
rect 1106 45616 1582 45684
rect 1106 45560 1130 45616
rect 1186 45560 1254 45616
rect 1310 45560 1378 45616
rect 1434 45560 1502 45616
rect 1558 45560 1582 45616
rect 1106 45492 1582 45560
rect 1106 45436 1130 45492
rect 1186 45436 1254 45492
rect 1310 45436 1378 45492
rect 1434 45436 1502 45492
rect 1558 45436 1582 45492
rect 1106 45424 1582 45436
rect 85788 45864 86264 45876
rect 85788 45808 85812 45864
rect 85868 45808 85936 45864
rect 85992 45808 86060 45864
rect 86116 45808 86184 45864
rect 86240 45808 86264 45864
rect 85788 45740 86264 45808
rect 85788 45684 85812 45740
rect 85868 45684 85936 45740
rect 85992 45684 86060 45740
rect 86116 45684 86184 45740
rect 86240 45684 86264 45740
rect 85788 45616 86264 45684
rect 85788 45560 85812 45616
rect 85868 45560 85936 45616
rect 85992 45560 86060 45616
rect 86116 45560 86184 45616
rect 86240 45560 86264 45616
rect 85788 45492 86264 45560
rect 85788 45436 85812 45492
rect 85868 45436 85936 45492
rect 85992 45436 86060 45492
rect 86116 45436 86184 45492
rect 86240 45436 86264 45492
rect 85788 45424 86264 45436
rect 86588 44964 87064 44976
rect 86588 44908 86612 44964
rect 86668 44908 86736 44964
rect 86792 44908 86860 44964
rect 86916 44908 86984 44964
rect 87040 44908 87064 44964
rect 1906 44840 2382 44900
rect 1906 44784 1930 44840
rect 1986 44784 2054 44840
rect 2110 44784 2178 44840
rect 2234 44784 2302 44840
rect 2358 44784 2382 44840
rect 1906 44716 2382 44784
rect 1906 44660 1930 44716
rect 1986 44660 2054 44716
rect 2110 44660 2178 44716
rect 2234 44660 2302 44716
rect 2358 44660 2382 44716
rect 1906 44600 2382 44660
rect 86588 44840 87064 44908
rect 86588 44784 86612 44840
rect 86668 44784 86736 44840
rect 86792 44784 86860 44840
rect 86916 44784 86984 44840
rect 87040 44784 87064 44840
rect 86588 44716 87064 44784
rect 86588 44660 86612 44716
rect 86668 44660 86736 44716
rect 86792 44660 86860 44716
rect 86916 44660 86984 44716
rect 87040 44660 87064 44716
rect 86588 44592 87064 44660
rect 86588 44536 86612 44592
rect 86668 44536 86736 44592
rect 86792 44536 86860 44592
rect 86916 44536 86984 44592
rect 87040 44536 87064 44592
rect 86588 44524 87064 44536
rect 1106 44064 1582 44076
rect 1106 44008 1130 44064
rect 1186 44008 1254 44064
rect 1310 44008 1378 44064
rect 1434 44008 1502 44064
rect 1558 44008 1582 44064
rect 1106 43940 1582 44008
rect 1106 43884 1130 43940
rect 1186 43884 1254 43940
rect 1310 43884 1378 43940
rect 1434 43884 1502 43940
rect 1558 43884 1582 43940
rect 1106 43816 1582 43884
rect 1106 43760 1130 43816
rect 1186 43760 1254 43816
rect 1310 43760 1378 43816
rect 1434 43760 1502 43816
rect 1558 43760 1582 43816
rect 1106 43692 1582 43760
rect 1106 43636 1130 43692
rect 1186 43636 1254 43692
rect 1310 43636 1378 43692
rect 1434 43636 1502 43692
rect 1558 43636 1582 43692
rect 1106 43624 1582 43636
rect 85788 44064 86264 44076
rect 85788 44008 85812 44064
rect 85868 44008 85936 44064
rect 85992 44008 86060 44064
rect 86116 44008 86184 44064
rect 86240 44008 86264 44064
rect 85788 43940 86264 44008
rect 85788 43884 85812 43940
rect 85868 43884 85936 43940
rect 85992 43884 86060 43940
rect 86116 43884 86184 43940
rect 86240 43884 86264 43940
rect 85788 43816 86264 43884
rect 85788 43760 85812 43816
rect 85868 43760 85936 43816
rect 85992 43760 86060 43816
rect 86116 43760 86184 43816
rect 86240 43760 86264 43816
rect 85788 43692 86264 43760
rect 85788 43636 85812 43692
rect 85868 43636 85936 43692
rect 85992 43636 86060 43692
rect 86116 43636 86184 43692
rect 86240 43636 86264 43692
rect 85788 43624 86264 43636
rect 86588 43164 87064 43176
rect 86588 43108 86612 43164
rect 86668 43108 86736 43164
rect 86792 43108 86860 43164
rect 86916 43108 86984 43164
rect 87040 43108 87064 43164
rect 1906 43040 2382 43100
rect 1906 42984 1930 43040
rect 1986 42984 2054 43040
rect 2110 42984 2178 43040
rect 2234 42984 2302 43040
rect 2358 42984 2382 43040
rect 1906 42916 2382 42984
rect 1906 42860 1930 42916
rect 1986 42860 2054 42916
rect 2110 42860 2178 42916
rect 2234 42860 2302 42916
rect 2358 42860 2382 42916
rect 1906 42800 2382 42860
rect 86588 43040 87064 43108
rect 86588 42984 86612 43040
rect 86668 42984 86736 43040
rect 86792 42984 86860 43040
rect 86916 42984 86984 43040
rect 87040 42984 87064 43040
rect 86588 42916 87064 42984
rect 86588 42860 86612 42916
rect 86668 42860 86736 42916
rect 86792 42860 86860 42916
rect 86916 42860 86984 42916
rect 87040 42860 87064 42916
rect 86588 42792 87064 42860
rect 86588 42736 86612 42792
rect 86668 42736 86736 42792
rect 86792 42736 86860 42792
rect 86916 42736 86984 42792
rect 87040 42736 87064 42792
rect 86588 42724 87064 42736
rect 1106 42264 1582 42276
rect 1106 42208 1130 42264
rect 1186 42208 1254 42264
rect 1310 42208 1378 42264
rect 1434 42208 1502 42264
rect 1558 42208 1582 42264
rect 1106 42140 1582 42208
rect 1106 42084 1130 42140
rect 1186 42084 1254 42140
rect 1310 42084 1378 42140
rect 1434 42084 1502 42140
rect 1558 42084 1582 42140
rect 1106 42016 1582 42084
rect 1106 41960 1130 42016
rect 1186 41960 1254 42016
rect 1310 41960 1378 42016
rect 1434 41960 1502 42016
rect 1558 41960 1582 42016
rect 1106 41892 1582 41960
rect 1106 41836 1130 41892
rect 1186 41836 1254 41892
rect 1310 41836 1378 41892
rect 1434 41836 1502 41892
rect 1558 41836 1582 41892
rect 1106 41824 1582 41836
rect 85788 42264 86264 42276
rect 85788 42208 85812 42264
rect 85868 42208 85936 42264
rect 85992 42208 86060 42264
rect 86116 42208 86184 42264
rect 86240 42208 86264 42264
rect 85788 42140 86264 42208
rect 85788 42084 85812 42140
rect 85868 42084 85936 42140
rect 85992 42084 86060 42140
rect 86116 42084 86184 42140
rect 86240 42084 86264 42140
rect 85788 42016 86264 42084
rect 85788 41960 85812 42016
rect 85868 41960 85936 42016
rect 85992 41960 86060 42016
rect 86116 41960 86184 42016
rect 86240 41960 86264 42016
rect 85788 41892 86264 41960
rect 85788 41836 85812 41892
rect 85868 41836 85936 41892
rect 85992 41836 86060 41892
rect 86116 41836 86184 41892
rect 86240 41836 86264 41892
rect 85788 41824 86264 41836
rect 86588 41364 87064 41376
rect 86588 41308 86612 41364
rect 86668 41308 86736 41364
rect 86792 41308 86860 41364
rect 86916 41308 86984 41364
rect 87040 41308 87064 41364
rect 1906 41240 2382 41300
rect 1906 41184 1930 41240
rect 1986 41184 2054 41240
rect 2110 41184 2178 41240
rect 2234 41184 2302 41240
rect 2358 41184 2382 41240
rect 1906 41116 2382 41184
rect 1906 41060 1930 41116
rect 1986 41060 2054 41116
rect 2110 41060 2178 41116
rect 2234 41060 2302 41116
rect 2358 41060 2382 41116
rect 1906 41000 2382 41060
rect 86588 41240 87064 41308
rect 86588 41184 86612 41240
rect 86668 41184 86736 41240
rect 86792 41184 86860 41240
rect 86916 41184 86984 41240
rect 87040 41184 87064 41240
rect 86588 41116 87064 41184
rect 86588 41060 86612 41116
rect 86668 41060 86736 41116
rect 86792 41060 86860 41116
rect 86916 41060 86984 41116
rect 87040 41060 87064 41116
rect 86588 40992 87064 41060
rect 86588 40936 86612 40992
rect 86668 40936 86736 40992
rect 86792 40936 86860 40992
rect 86916 40936 86984 40992
rect 87040 40936 87064 40992
rect 86588 40924 87064 40936
rect 1106 40464 1582 40476
rect 1106 40408 1130 40464
rect 1186 40408 1254 40464
rect 1310 40408 1378 40464
rect 1434 40408 1502 40464
rect 1558 40408 1582 40464
rect 1106 40340 1582 40408
rect 1106 40284 1130 40340
rect 1186 40284 1254 40340
rect 1310 40284 1378 40340
rect 1434 40284 1502 40340
rect 1558 40284 1582 40340
rect 1106 40216 1582 40284
rect 1106 40160 1130 40216
rect 1186 40160 1254 40216
rect 1310 40160 1378 40216
rect 1434 40160 1502 40216
rect 1558 40160 1582 40216
rect 1106 40092 1582 40160
rect 1106 40036 1130 40092
rect 1186 40036 1254 40092
rect 1310 40036 1378 40092
rect 1434 40036 1502 40092
rect 1558 40036 1582 40092
rect 1106 40024 1582 40036
rect 85788 40464 86264 40476
rect 85788 40408 85812 40464
rect 85868 40408 85936 40464
rect 85992 40408 86060 40464
rect 86116 40408 86184 40464
rect 86240 40408 86264 40464
rect 85788 40340 86264 40408
rect 85788 40284 85812 40340
rect 85868 40284 85936 40340
rect 85992 40284 86060 40340
rect 86116 40284 86184 40340
rect 86240 40284 86264 40340
rect 85788 40216 86264 40284
rect 85788 40160 85812 40216
rect 85868 40160 85936 40216
rect 85992 40160 86060 40216
rect 86116 40160 86184 40216
rect 86240 40160 86264 40216
rect 85788 40092 86264 40160
rect 85788 40036 85812 40092
rect 85868 40036 85936 40092
rect 85992 40036 86060 40092
rect 86116 40036 86184 40092
rect 86240 40036 86264 40092
rect 85788 40024 86264 40036
rect 86588 39564 87064 39576
rect 86588 39508 86612 39564
rect 86668 39508 86736 39564
rect 86792 39508 86860 39564
rect 86916 39508 86984 39564
rect 87040 39508 87064 39564
rect 1906 39440 2382 39500
rect 1906 39384 1930 39440
rect 1986 39384 2054 39440
rect 2110 39384 2178 39440
rect 2234 39384 2302 39440
rect 2358 39384 2382 39440
rect 1906 39316 2382 39384
rect 1906 39260 1930 39316
rect 1986 39260 2054 39316
rect 2110 39260 2178 39316
rect 2234 39260 2302 39316
rect 2358 39260 2382 39316
rect 1906 39200 2382 39260
rect 86588 39440 87064 39508
rect 86588 39384 86612 39440
rect 86668 39384 86736 39440
rect 86792 39384 86860 39440
rect 86916 39384 86984 39440
rect 87040 39384 87064 39440
rect 86588 39316 87064 39384
rect 86588 39260 86612 39316
rect 86668 39260 86736 39316
rect 86792 39260 86860 39316
rect 86916 39260 86984 39316
rect 87040 39260 87064 39316
rect 86588 39192 87064 39260
rect 86588 39136 86612 39192
rect 86668 39136 86736 39192
rect 86792 39136 86860 39192
rect 86916 39136 86984 39192
rect 87040 39136 87064 39192
rect 86588 39124 87064 39136
rect 1106 38664 1582 38676
rect 1106 38608 1130 38664
rect 1186 38608 1254 38664
rect 1310 38608 1378 38664
rect 1434 38608 1502 38664
rect 1558 38608 1582 38664
rect 1106 38540 1582 38608
rect 1106 38484 1130 38540
rect 1186 38484 1254 38540
rect 1310 38484 1378 38540
rect 1434 38484 1502 38540
rect 1558 38484 1582 38540
rect 1106 38416 1582 38484
rect 1106 38360 1130 38416
rect 1186 38360 1254 38416
rect 1310 38360 1378 38416
rect 1434 38360 1502 38416
rect 1558 38360 1582 38416
rect 1106 38292 1582 38360
rect 1106 38236 1130 38292
rect 1186 38236 1254 38292
rect 1310 38236 1378 38292
rect 1434 38236 1502 38292
rect 1558 38236 1582 38292
rect 1106 38224 1582 38236
rect 85788 38664 86264 38676
rect 85788 38608 85812 38664
rect 85868 38608 85936 38664
rect 85992 38608 86060 38664
rect 86116 38608 86184 38664
rect 86240 38608 86264 38664
rect 85788 38540 86264 38608
rect 85788 38484 85812 38540
rect 85868 38484 85936 38540
rect 85992 38484 86060 38540
rect 86116 38484 86184 38540
rect 86240 38484 86264 38540
rect 85788 38416 86264 38484
rect 85788 38360 85812 38416
rect 85868 38360 85936 38416
rect 85992 38360 86060 38416
rect 86116 38360 86184 38416
rect 86240 38360 86264 38416
rect 85788 38292 86264 38360
rect 85788 38236 85812 38292
rect 85868 38236 85936 38292
rect 85992 38236 86060 38292
rect 86116 38236 86184 38292
rect 86240 38236 86264 38292
rect 85788 38224 86264 38236
rect 86588 37764 87064 37776
rect 86588 37708 86612 37764
rect 86668 37708 86736 37764
rect 86792 37708 86860 37764
rect 86916 37708 86984 37764
rect 87040 37708 87064 37764
rect 1906 37640 2382 37700
rect 1906 37584 1930 37640
rect 1986 37584 2054 37640
rect 2110 37584 2178 37640
rect 2234 37584 2302 37640
rect 2358 37584 2382 37640
rect 1906 37516 2382 37584
rect 1906 37460 1930 37516
rect 1986 37460 2054 37516
rect 2110 37460 2178 37516
rect 2234 37460 2302 37516
rect 2358 37460 2382 37516
rect 1906 37400 2382 37460
rect 86588 37640 87064 37708
rect 86588 37584 86612 37640
rect 86668 37584 86736 37640
rect 86792 37584 86860 37640
rect 86916 37584 86984 37640
rect 87040 37584 87064 37640
rect 86588 37516 87064 37584
rect 86588 37460 86612 37516
rect 86668 37460 86736 37516
rect 86792 37460 86860 37516
rect 86916 37460 86984 37516
rect 87040 37460 87064 37516
rect 86588 37392 87064 37460
rect 86588 37336 86612 37392
rect 86668 37336 86736 37392
rect 86792 37336 86860 37392
rect 86916 37336 86984 37392
rect 87040 37336 87064 37392
rect 86588 37324 87064 37336
rect 1106 36864 1582 36876
rect 1106 36808 1130 36864
rect 1186 36808 1254 36864
rect 1310 36808 1378 36864
rect 1434 36808 1502 36864
rect 1558 36808 1582 36864
rect 1106 36740 1582 36808
rect 1106 36684 1130 36740
rect 1186 36684 1254 36740
rect 1310 36684 1378 36740
rect 1434 36684 1502 36740
rect 1558 36684 1582 36740
rect 1106 36616 1582 36684
rect 1106 36560 1130 36616
rect 1186 36560 1254 36616
rect 1310 36560 1378 36616
rect 1434 36560 1502 36616
rect 1558 36560 1582 36616
rect 1106 36492 1582 36560
rect 1106 36436 1130 36492
rect 1186 36436 1254 36492
rect 1310 36436 1378 36492
rect 1434 36436 1502 36492
rect 1558 36436 1582 36492
rect 1106 36424 1582 36436
rect 85788 36864 86264 36876
rect 85788 36808 85812 36864
rect 85868 36808 85936 36864
rect 85992 36808 86060 36864
rect 86116 36808 86184 36864
rect 86240 36808 86264 36864
rect 85788 36740 86264 36808
rect 85788 36684 85812 36740
rect 85868 36684 85936 36740
rect 85992 36684 86060 36740
rect 86116 36684 86184 36740
rect 86240 36684 86264 36740
rect 85788 36616 86264 36684
rect 85788 36560 85812 36616
rect 85868 36560 85936 36616
rect 85992 36560 86060 36616
rect 86116 36560 86184 36616
rect 86240 36560 86264 36616
rect 85788 36492 86264 36560
rect 85788 36436 85812 36492
rect 85868 36436 85936 36492
rect 85992 36436 86060 36492
rect 86116 36436 86184 36492
rect 86240 36436 86264 36492
rect 85788 36424 86264 36436
rect 86588 35964 87064 35976
rect 86588 35908 86612 35964
rect 86668 35908 86736 35964
rect 86792 35908 86860 35964
rect 86916 35908 86984 35964
rect 87040 35908 87064 35964
rect 1906 35840 2382 35900
rect 1906 35784 1930 35840
rect 1986 35784 2054 35840
rect 2110 35784 2178 35840
rect 2234 35784 2302 35840
rect 2358 35784 2382 35840
rect 1906 35716 2382 35784
rect 1906 35660 1930 35716
rect 1986 35660 2054 35716
rect 2110 35660 2178 35716
rect 2234 35660 2302 35716
rect 2358 35660 2382 35716
rect 1906 35600 2382 35660
rect 86588 35840 87064 35908
rect 86588 35784 86612 35840
rect 86668 35784 86736 35840
rect 86792 35784 86860 35840
rect 86916 35784 86984 35840
rect 87040 35784 87064 35840
rect 86588 35716 87064 35784
rect 86588 35660 86612 35716
rect 86668 35660 86736 35716
rect 86792 35660 86860 35716
rect 86916 35660 86984 35716
rect 87040 35660 87064 35716
rect 86588 35592 87064 35660
rect 86588 35536 86612 35592
rect 86668 35536 86736 35592
rect 86792 35536 86860 35592
rect 86916 35536 86984 35592
rect 87040 35536 87064 35592
rect 86588 35524 87064 35536
rect 1106 35064 1582 35076
rect 1106 35008 1130 35064
rect 1186 35008 1254 35064
rect 1310 35008 1378 35064
rect 1434 35008 1502 35064
rect 1558 35008 1582 35064
rect 1106 34940 1582 35008
rect 1106 34884 1130 34940
rect 1186 34884 1254 34940
rect 1310 34884 1378 34940
rect 1434 34884 1502 34940
rect 1558 34884 1582 34940
rect 1106 34816 1582 34884
rect 1106 34760 1130 34816
rect 1186 34760 1254 34816
rect 1310 34760 1378 34816
rect 1434 34760 1502 34816
rect 1558 34760 1582 34816
rect 1106 34692 1582 34760
rect 1106 34636 1130 34692
rect 1186 34636 1254 34692
rect 1310 34636 1378 34692
rect 1434 34636 1502 34692
rect 1558 34636 1582 34692
rect 1106 34624 1582 34636
rect 85788 35064 86264 35076
rect 85788 35008 85812 35064
rect 85868 35008 85936 35064
rect 85992 35008 86060 35064
rect 86116 35008 86184 35064
rect 86240 35008 86264 35064
rect 85788 34940 86264 35008
rect 85788 34884 85812 34940
rect 85868 34884 85936 34940
rect 85992 34884 86060 34940
rect 86116 34884 86184 34940
rect 86240 34884 86264 34940
rect 85788 34816 86264 34884
rect 85788 34760 85812 34816
rect 85868 34760 85936 34816
rect 85992 34760 86060 34816
rect 86116 34760 86184 34816
rect 86240 34760 86264 34816
rect 85788 34692 86264 34760
rect 85788 34636 85812 34692
rect 85868 34636 85936 34692
rect 85992 34636 86060 34692
rect 86116 34636 86184 34692
rect 86240 34636 86264 34692
rect 85788 34624 86264 34636
rect 86588 34164 87064 34176
rect 86588 34108 86612 34164
rect 86668 34108 86736 34164
rect 86792 34108 86860 34164
rect 86916 34108 86984 34164
rect 87040 34108 87064 34164
rect 1906 34040 2382 34100
rect 1906 33984 1930 34040
rect 1986 33984 2054 34040
rect 2110 33984 2178 34040
rect 2234 33984 2302 34040
rect 2358 33984 2382 34040
rect 1906 33916 2382 33984
rect 1906 33860 1930 33916
rect 1986 33860 2054 33916
rect 2110 33860 2178 33916
rect 2234 33860 2302 33916
rect 2358 33860 2382 33916
rect 1906 33800 2382 33860
rect 86588 34040 87064 34108
rect 86588 33984 86612 34040
rect 86668 33984 86736 34040
rect 86792 33984 86860 34040
rect 86916 33984 86984 34040
rect 87040 33984 87064 34040
rect 86588 33916 87064 33984
rect 86588 33860 86612 33916
rect 86668 33860 86736 33916
rect 86792 33860 86860 33916
rect 86916 33860 86984 33916
rect 87040 33860 87064 33916
rect 86588 33792 87064 33860
rect 86588 33736 86612 33792
rect 86668 33736 86736 33792
rect 86792 33736 86860 33792
rect 86916 33736 86984 33792
rect 87040 33736 87064 33792
rect 86588 33724 87064 33736
rect 1106 33264 1582 33276
rect 1106 33208 1130 33264
rect 1186 33208 1254 33264
rect 1310 33208 1378 33264
rect 1434 33208 1502 33264
rect 1558 33208 1582 33264
rect 1106 33140 1582 33208
rect 1106 33084 1130 33140
rect 1186 33084 1254 33140
rect 1310 33084 1378 33140
rect 1434 33084 1502 33140
rect 1558 33084 1582 33140
rect 1106 33016 1582 33084
rect 1106 32960 1130 33016
rect 1186 32960 1254 33016
rect 1310 32960 1378 33016
rect 1434 32960 1502 33016
rect 1558 32960 1582 33016
rect 1106 32892 1582 32960
rect 1106 32836 1130 32892
rect 1186 32836 1254 32892
rect 1310 32836 1378 32892
rect 1434 32836 1502 32892
rect 1558 32836 1582 32892
rect 1106 32824 1582 32836
rect 85788 33264 86264 33276
rect 85788 33208 85812 33264
rect 85868 33208 85936 33264
rect 85992 33208 86060 33264
rect 86116 33208 86184 33264
rect 86240 33208 86264 33264
rect 85788 33140 86264 33208
rect 85788 33084 85812 33140
rect 85868 33084 85936 33140
rect 85992 33084 86060 33140
rect 86116 33084 86184 33140
rect 86240 33084 86264 33140
rect 85788 33016 86264 33084
rect 85788 32960 85812 33016
rect 85868 32960 85936 33016
rect 85992 32960 86060 33016
rect 86116 32960 86184 33016
rect 86240 32960 86264 33016
rect 85788 32892 86264 32960
rect 85788 32836 85812 32892
rect 85868 32836 85936 32892
rect 85992 32836 86060 32892
rect 86116 32836 86184 32892
rect 86240 32836 86264 32892
rect 85788 32824 86264 32836
rect 86588 32364 87064 32376
rect 86588 32308 86612 32364
rect 86668 32308 86736 32364
rect 86792 32308 86860 32364
rect 86916 32308 86984 32364
rect 87040 32308 87064 32364
rect 1906 32240 2382 32300
rect 1906 32184 1930 32240
rect 1986 32184 2054 32240
rect 2110 32184 2178 32240
rect 2234 32184 2302 32240
rect 2358 32184 2382 32240
rect 1906 32116 2382 32184
rect 1906 32060 1930 32116
rect 1986 32060 2054 32116
rect 2110 32060 2178 32116
rect 2234 32060 2302 32116
rect 2358 32060 2382 32116
rect 1906 32000 2382 32060
rect 86588 32240 87064 32308
rect 86588 32184 86612 32240
rect 86668 32184 86736 32240
rect 86792 32184 86860 32240
rect 86916 32184 86984 32240
rect 87040 32184 87064 32240
rect 86588 32116 87064 32184
rect 86588 32060 86612 32116
rect 86668 32060 86736 32116
rect 86792 32060 86860 32116
rect 86916 32060 86984 32116
rect 87040 32060 87064 32116
rect 86588 31992 87064 32060
rect 86588 31936 86612 31992
rect 86668 31936 86736 31992
rect 86792 31936 86860 31992
rect 86916 31936 86984 31992
rect 87040 31936 87064 31992
rect 86588 31924 87064 31936
rect 1106 31464 1582 31476
rect 1106 31408 1130 31464
rect 1186 31408 1254 31464
rect 1310 31408 1378 31464
rect 1434 31408 1502 31464
rect 1558 31408 1582 31464
rect 1106 31340 1582 31408
rect 1106 31284 1130 31340
rect 1186 31284 1254 31340
rect 1310 31284 1378 31340
rect 1434 31284 1502 31340
rect 1558 31284 1582 31340
rect 1106 31216 1582 31284
rect 1106 31160 1130 31216
rect 1186 31160 1254 31216
rect 1310 31160 1378 31216
rect 1434 31160 1502 31216
rect 1558 31160 1582 31216
rect 1106 31092 1582 31160
rect 1106 31036 1130 31092
rect 1186 31036 1254 31092
rect 1310 31036 1378 31092
rect 1434 31036 1502 31092
rect 1558 31036 1582 31092
rect 1106 31024 1582 31036
rect 85788 31464 86264 31476
rect 85788 31408 85812 31464
rect 85868 31408 85936 31464
rect 85992 31408 86060 31464
rect 86116 31408 86184 31464
rect 86240 31408 86264 31464
rect 85788 31340 86264 31408
rect 85788 31284 85812 31340
rect 85868 31284 85936 31340
rect 85992 31284 86060 31340
rect 86116 31284 86184 31340
rect 86240 31284 86264 31340
rect 85788 31216 86264 31284
rect 85788 31160 85812 31216
rect 85868 31160 85936 31216
rect 85992 31160 86060 31216
rect 86116 31160 86184 31216
rect 86240 31160 86264 31216
rect 85788 31092 86264 31160
rect 85788 31036 85812 31092
rect 85868 31036 85936 31092
rect 85992 31036 86060 31092
rect 86116 31036 86184 31092
rect 86240 31036 86264 31092
rect 85788 31024 86264 31036
rect 86588 30564 87064 30576
rect 86588 30508 86612 30564
rect 86668 30508 86736 30564
rect 86792 30508 86860 30564
rect 86916 30508 86984 30564
rect 87040 30508 87064 30564
rect 1906 30440 2382 30500
rect 1906 30384 1930 30440
rect 1986 30384 2054 30440
rect 2110 30384 2178 30440
rect 2234 30384 2302 30440
rect 2358 30384 2382 30440
rect 1906 30316 2382 30384
rect 1906 30260 1930 30316
rect 1986 30260 2054 30316
rect 2110 30260 2178 30316
rect 2234 30260 2302 30316
rect 2358 30260 2382 30316
rect 1906 30200 2382 30260
rect 86588 30440 87064 30508
rect 86588 30384 86612 30440
rect 86668 30384 86736 30440
rect 86792 30384 86860 30440
rect 86916 30384 86984 30440
rect 87040 30384 87064 30440
rect 86588 30316 87064 30384
rect 86588 30260 86612 30316
rect 86668 30260 86736 30316
rect 86792 30260 86860 30316
rect 86916 30260 86984 30316
rect 87040 30260 87064 30316
rect 86588 30192 87064 30260
rect 86588 30136 86612 30192
rect 86668 30136 86736 30192
rect 86792 30136 86860 30192
rect 86916 30136 86984 30192
rect 87040 30136 87064 30192
rect 86588 30124 87064 30136
rect 1106 29664 1582 29676
rect 1106 29608 1130 29664
rect 1186 29608 1254 29664
rect 1310 29608 1378 29664
rect 1434 29608 1502 29664
rect 1558 29608 1582 29664
rect 1106 29540 1582 29608
rect 1106 29484 1130 29540
rect 1186 29484 1254 29540
rect 1310 29484 1378 29540
rect 1434 29484 1502 29540
rect 1558 29484 1582 29540
rect 1106 29416 1582 29484
rect 1106 29360 1130 29416
rect 1186 29360 1254 29416
rect 1310 29360 1378 29416
rect 1434 29360 1502 29416
rect 1558 29360 1582 29416
rect 1106 29292 1582 29360
rect 1106 29236 1130 29292
rect 1186 29236 1254 29292
rect 1310 29236 1378 29292
rect 1434 29236 1502 29292
rect 1558 29236 1582 29292
rect 1106 29224 1582 29236
rect 85788 29664 86264 29676
rect 85788 29608 85812 29664
rect 85868 29608 85936 29664
rect 85992 29608 86060 29664
rect 86116 29608 86184 29664
rect 86240 29608 86264 29664
rect 85788 29540 86264 29608
rect 85788 29484 85812 29540
rect 85868 29484 85936 29540
rect 85992 29484 86060 29540
rect 86116 29484 86184 29540
rect 86240 29484 86264 29540
rect 85788 29416 86264 29484
rect 85788 29360 85812 29416
rect 85868 29360 85936 29416
rect 85992 29360 86060 29416
rect 86116 29360 86184 29416
rect 86240 29360 86264 29416
rect 85788 29292 86264 29360
rect 85788 29236 85812 29292
rect 85868 29236 85936 29292
rect 85992 29236 86060 29292
rect 86116 29236 86184 29292
rect 86240 29236 86264 29292
rect 85788 29224 86264 29236
rect 86588 28764 87064 28776
rect 86588 28708 86612 28764
rect 86668 28708 86736 28764
rect 86792 28708 86860 28764
rect 86916 28708 86984 28764
rect 87040 28708 87064 28764
rect 1906 28640 2382 28700
rect 1906 28584 1930 28640
rect 1986 28584 2054 28640
rect 2110 28584 2178 28640
rect 2234 28584 2302 28640
rect 2358 28584 2382 28640
rect 1906 28516 2382 28584
rect 1906 28460 1930 28516
rect 1986 28460 2054 28516
rect 2110 28460 2178 28516
rect 2234 28460 2302 28516
rect 2358 28460 2382 28516
rect 1906 28400 2382 28460
rect 86588 28640 87064 28708
rect 86588 28584 86612 28640
rect 86668 28584 86736 28640
rect 86792 28584 86860 28640
rect 86916 28584 86984 28640
rect 87040 28584 87064 28640
rect 86588 28516 87064 28584
rect 86588 28460 86612 28516
rect 86668 28460 86736 28516
rect 86792 28460 86860 28516
rect 86916 28460 86984 28516
rect 87040 28460 87064 28516
rect 86588 28392 87064 28460
rect 86588 28336 86612 28392
rect 86668 28336 86736 28392
rect 86792 28336 86860 28392
rect 86916 28336 86984 28392
rect 87040 28336 87064 28392
rect 86588 28324 87064 28336
rect 1106 27864 1582 27876
rect 1106 27808 1130 27864
rect 1186 27808 1254 27864
rect 1310 27808 1378 27864
rect 1434 27808 1502 27864
rect 1558 27808 1582 27864
rect 1106 27740 1582 27808
rect 1106 27684 1130 27740
rect 1186 27684 1254 27740
rect 1310 27684 1378 27740
rect 1434 27684 1502 27740
rect 1558 27684 1582 27740
rect 1106 27616 1582 27684
rect 1106 27560 1130 27616
rect 1186 27560 1254 27616
rect 1310 27560 1378 27616
rect 1434 27560 1502 27616
rect 1558 27560 1582 27616
rect 1106 27492 1582 27560
rect 1106 27436 1130 27492
rect 1186 27436 1254 27492
rect 1310 27436 1378 27492
rect 1434 27436 1502 27492
rect 1558 27436 1582 27492
rect 1106 27424 1582 27436
rect 85788 27864 86264 27876
rect 85788 27808 85812 27864
rect 85868 27808 85936 27864
rect 85992 27808 86060 27864
rect 86116 27808 86184 27864
rect 86240 27808 86264 27864
rect 85788 27740 86264 27808
rect 85788 27684 85812 27740
rect 85868 27684 85936 27740
rect 85992 27684 86060 27740
rect 86116 27684 86184 27740
rect 86240 27684 86264 27740
rect 85788 27616 86264 27684
rect 85788 27560 85812 27616
rect 85868 27560 85936 27616
rect 85992 27560 86060 27616
rect 86116 27560 86184 27616
rect 86240 27560 86264 27616
rect 85788 27492 86264 27560
rect 85788 27436 85812 27492
rect 85868 27436 85936 27492
rect 85992 27436 86060 27492
rect 86116 27436 86184 27492
rect 86240 27436 86264 27492
rect 85788 27424 86264 27436
rect 86588 26964 87064 26976
rect 86588 26908 86612 26964
rect 86668 26908 86736 26964
rect 86792 26908 86860 26964
rect 86916 26908 86984 26964
rect 87040 26908 87064 26964
rect 1906 26840 2382 26900
rect 1906 26784 1930 26840
rect 1986 26784 2054 26840
rect 2110 26784 2178 26840
rect 2234 26784 2302 26840
rect 2358 26784 2382 26840
rect 1906 26716 2382 26784
rect 1906 26660 1930 26716
rect 1986 26660 2054 26716
rect 2110 26660 2178 26716
rect 2234 26660 2302 26716
rect 2358 26660 2382 26716
rect 1906 26600 2382 26660
rect 86588 26840 87064 26908
rect 86588 26784 86612 26840
rect 86668 26784 86736 26840
rect 86792 26784 86860 26840
rect 86916 26784 86984 26840
rect 87040 26784 87064 26840
rect 86588 26716 87064 26784
rect 86588 26660 86612 26716
rect 86668 26660 86736 26716
rect 86792 26660 86860 26716
rect 86916 26660 86984 26716
rect 87040 26660 87064 26716
rect 86588 26592 87064 26660
rect 86588 26536 86612 26592
rect 86668 26536 86736 26592
rect 86792 26536 86860 26592
rect 86916 26536 86984 26592
rect 87040 26536 87064 26592
rect 86588 26524 87064 26536
rect 1106 26064 1582 26076
rect 1106 26008 1130 26064
rect 1186 26008 1254 26064
rect 1310 26008 1378 26064
rect 1434 26008 1502 26064
rect 1558 26008 1582 26064
rect 1106 25940 1582 26008
rect 1106 25884 1130 25940
rect 1186 25884 1254 25940
rect 1310 25884 1378 25940
rect 1434 25884 1502 25940
rect 1558 25884 1582 25940
rect 1106 25816 1582 25884
rect 1106 25760 1130 25816
rect 1186 25760 1254 25816
rect 1310 25760 1378 25816
rect 1434 25760 1502 25816
rect 1558 25760 1582 25816
rect 1106 25692 1582 25760
rect 1106 25636 1130 25692
rect 1186 25636 1254 25692
rect 1310 25636 1378 25692
rect 1434 25636 1502 25692
rect 1558 25636 1582 25692
rect 1106 25624 1582 25636
rect 85788 26064 86264 26076
rect 85788 26008 85812 26064
rect 85868 26008 85936 26064
rect 85992 26008 86060 26064
rect 86116 26008 86184 26064
rect 86240 26008 86264 26064
rect 85788 25940 86264 26008
rect 85788 25884 85812 25940
rect 85868 25884 85936 25940
rect 85992 25884 86060 25940
rect 86116 25884 86184 25940
rect 86240 25884 86264 25940
rect 85788 25816 86264 25884
rect 85788 25760 85812 25816
rect 85868 25760 85936 25816
rect 85992 25760 86060 25816
rect 86116 25760 86184 25816
rect 86240 25760 86264 25816
rect 85788 25692 86264 25760
rect 85788 25636 85812 25692
rect 85868 25636 85936 25692
rect 85992 25636 86060 25692
rect 86116 25636 86184 25692
rect 86240 25636 86264 25692
rect 85788 25624 86264 25636
rect 86588 25164 87064 25176
rect 86588 25108 86612 25164
rect 86668 25108 86736 25164
rect 86792 25108 86860 25164
rect 86916 25108 86984 25164
rect 87040 25108 87064 25164
rect 1906 25040 2382 25100
rect 1906 24984 1930 25040
rect 1986 24984 2054 25040
rect 2110 24984 2178 25040
rect 2234 24984 2302 25040
rect 2358 24984 2382 25040
rect 1906 24916 2382 24984
rect 1906 24860 1930 24916
rect 1986 24860 2054 24916
rect 2110 24860 2178 24916
rect 2234 24860 2302 24916
rect 2358 24860 2382 24916
rect 1906 24800 2382 24860
rect 86588 25040 87064 25108
rect 86588 24984 86612 25040
rect 86668 24984 86736 25040
rect 86792 24984 86860 25040
rect 86916 24984 86984 25040
rect 87040 24984 87064 25040
rect 86588 24916 87064 24984
rect 86588 24860 86612 24916
rect 86668 24860 86736 24916
rect 86792 24860 86860 24916
rect 86916 24860 86984 24916
rect 87040 24860 87064 24916
rect 86588 24792 87064 24860
rect 86588 24736 86612 24792
rect 86668 24736 86736 24792
rect 86792 24736 86860 24792
rect 86916 24736 86984 24792
rect 87040 24736 87064 24792
rect 86588 24724 87064 24736
rect 1106 24264 1582 24276
rect 1106 24208 1130 24264
rect 1186 24208 1254 24264
rect 1310 24208 1378 24264
rect 1434 24208 1502 24264
rect 1558 24208 1582 24264
rect 1106 24140 1582 24208
rect 1106 24084 1130 24140
rect 1186 24084 1254 24140
rect 1310 24084 1378 24140
rect 1434 24084 1502 24140
rect 1558 24084 1582 24140
rect 1106 24016 1582 24084
rect 1106 23960 1130 24016
rect 1186 23960 1254 24016
rect 1310 23960 1378 24016
rect 1434 23960 1502 24016
rect 1558 23960 1582 24016
rect 1106 23892 1582 23960
rect 1106 23836 1130 23892
rect 1186 23836 1254 23892
rect 1310 23836 1378 23892
rect 1434 23836 1502 23892
rect 1558 23836 1582 23892
rect 1106 23824 1582 23836
rect 85788 24264 86264 24276
rect 85788 24208 85812 24264
rect 85868 24208 85936 24264
rect 85992 24208 86060 24264
rect 86116 24208 86184 24264
rect 86240 24208 86264 24264
rect 85788 24140 86264 24208
rect 85788 24084 85812 24140
rect 85868 24084 85936 24140
rect 85992 24084 86060 24140
rect 86116 24084 86184 24140
rect 86240 24084 86264 24140
rect 85788 24016 86264 24084
rect 85788 23960 85812 24016
rect 85868 23960 85936 24016
rect 85992 23960 86060 24016
rect 86116 23960 86184 24016
rect 86240 23960 86264 24016
rect 85788 23892 86264 23960
rect 85788 23836 85812 23892
rect 85868 23836 85936 23892
rect 85992 23836 86060 23892
rect 86116 23836 86184 23892
rect 86240 23836 86264 23892
rect 85788 23824 86264 23836
rect 86588 23364 87064 23376
rect 86588 23308 86612 23364
rect 86668 23308 86736 23364
rect 86792 23308 86860 23364
rect 86916 23308 86984 23364
rect 87040 23308 87064 23364
rect 1906 23240 2382 23300
rect 1906 23184 1930 23240
rect 1986 23184 2054 23240
rect 2110 23184 2178 23240
rect 2234 23184 2302 23240
rect 2358 23184 2382 23240
rect 1906 23116 2382 23184
rect 1906 23060 1930 23116
rect 1986 23060 2054 23116
rect 2110 23060 2178 23116
rect 2234 23060 2302 23116
rect 2358 23060 2382 23116
rect 1906 23000 2382 23060
rect 86588 23240 87064 23308
rect 86588 23184 86612 23240
rect 86668 23184 86736 23240
rect 86792 23184 86860 23240
rect 86916 23184 86984 23240
rect 87040 23184 87064 23240
rect 86588 23116 87064 23184
rect 86588 23060 86612 23116
rect 86668 23060 86736 23116
rect 86792 23060 86860 23116
rect 86916 23060 86984 23116
rect 87040 23060 87064 23116
rect 86588 22992 87064 23060
rect 86588 22936 86612 22992
rect 86668 22936 86736 22992
rect 86792 22936 86860 22992
rect 86916 22936 86984 22992
rect 87040 22936 87064 22992
rect 86588 22924 87064 22936
rect 1106 22464 1582 22476
rect 1106 22408 1130 22464
rect 1186 22408 1254 22464
rect 1310 22408 1378 22464
rect 1434 22408 1502 22464
rect 1558 22408 1582 22464
rect 1106 22340 1582 22408
rect 1106 22284 1130 22340
rect 1186 22284 1254 22340
rect 1310 22284 1378 22340
rect 1434 22284 1502 22340
rect 1558 22284 1582 22340
rect 1106 22216 1582 22284
rect 1106 22160 1130 22216
rect 1186 22160 1254 22216
rect 1310 22160 1378 22216
rect 1434 22160 1502 22216
rect 1558 22160 1582 22216
rect 1106 22092 1582 22160
rect 1106 22036 1130 22092
rect 1186 22036 1254 22092
rect 1310 22036 1378 22092
rect 1434 22036 1502 22092
rect 1558 22036 1582 22092
rect 1106 22024 1582 22036
rect 85788 22464 86264 22476
rect 85788 22408 85812 22464
rect 85868 22408 85936 22464
rect 85992 22408 86060 22464
rect 86116 22408 86184 22464
rect 86240 22408 86264 22464
rect 85788 22340 86264 22408
rect 85788 22284 85812 22340
rect 85868 22284 85936 22340
rect 85992 22284 86060 22340
rect 86116 22284 86184 22340
rect 86240 22284 86264 22340
rect 85788 22216 86264 22284
rect 85788 22160 85812 22216
rect 85868 22160 85936 22216
rect 85992 22160 86060 22216
rect 86116 22160 86184 22216
rect 86240 22160 86264 22216
rect 85788 22092 86264 22160
rect 85788 22036 85812 22092
rect 85868 22036 85936 22092
rect 85992 22036 86060 22092
rect 86116 22036 86184 22092
rect 86240 22036 86264 22092
rect 85788 22024 86264 22036
rect 86588 21564 87064 21576
rect 86588 21508 86612 21564
rect 86668 21508 86736 21564
rect 86792 21508 86860 21564
rect 86916 21508 86984 21564
rect 87040 21508 87064 21564
rect 1906 21440 2382 21500
rect 1906 21384 1930 21440
rect 1986 21384 2054 21440
rect 2110 21384 2178 21440
rect 2234 21384 2302 21440
rect 2358 21384 2382 21440
rect 1906 21316 2382 21384
rect 1906 21260 1930 21316
rect 1986 21260 2054 21316
rect 2110 21260 2178 21316
rect 2234 21260 2302 21316
rect 2358 21260 2382 21316
rect 1906 21200 2382 21260
rect 86588 21440 87064 21508
rect 86588 21384 86612 21440
rect 86668 21384 86736 21440
rect 86792 21384 86860 21440
rect 86916 21384 86984 21440
rect 87040 21384 87064 21440
rect 86588 21316 87064 21384
rect 86588 21260 86612 21316
rect 86668 21260 86736 21316
rect 86792 21260 86860 21316
rect 86916 21260 86984 21316
rect 87040 21260 87064 21316
rect 86588 21192 87064 21260
rect 86588 21136 86612 21192
rect 86668 21136 86736 21192
rect 86792 21136 86860 21192
rect 86916 21136 86984 21192
rect 87040 21136 87064 21192
rect 86588 21124 87064 21136
rect 1106 20664 1582 20676
rect 1106 20608 1130 20664
rect 1186 20608 1254 20664
rect 1310 20608 1378 20664
rect 1434 20608 1502 20664
rect 1558 20608 1582 20664
rect 1106 20540 1582 20608
rect 1106 20484 1130 20540
rect 1186 20484 1254 20540
rect 1310 20484 1378 20540
rect 1434 20484 1502 20540
rect 1558 20484 1582 20540
rect 1106 20416 1582 20484
rect 1106 20360 1130 20416
rect 1186 20360 1254 20416
rect 1310 20360 1378 20416
rect 1434 20360 1502 20416
rect 1558 20360 1582 20416
rect 1106 20292 1582 20360
rect 1106 20236 1130 20292
rect 1186 20236 1254 20292
rect 1310 20236 1378 20292
rect 1434 20236 1502 20292
rect 1558 20236 1582 20292
rect 1106 20224 1582 20236
rect 85788 20664 86264 20676
rect 85788 20608 85812 20664
rect 85868 20608 85936 20664
rect 85992 20608 86060 20664
rect 86116 20608 86184 20664
rect 86240 20608 86264 20664
rect 85788 20540 86264 20608
rect 85788 20484 85812 20540
rect 85868 20484 85936 20540
rect 85992 20484 86060 20540
rect 86116 20484 86184 20540
rect 86240 20484 86264 20540
rect 85788 20416 86264 20484
rect 85788 20360 85812 20416
rect 85868 20360 85936 20416
rect 85992 20360 86060 20416
rect 86116 20360 86184 20416
rect 86240 20360 86264 20416
rect 85788 20292 86264 20360
rect 85788 20236 85812 20292
rect 85868 20236 85936 20292
rect 85992 20236 86060 20292
rect 86116 20236 86184 20292
rect 86240 20236 86264 20292
rect 85788 20224 86264 20236
rect 86588 19764 87064 19776
rect 86588 19708 86612 19764
rect 86668 19708 86736 19764
rect 86792 19708 86860 19764
rect 86916 19708 86984 19764
rect 87040 19708 87064 19764
rect 1906 19640 2382 19700
rect 1906 19584 1930 19640
rect 1986 19584 2054 19640
rect 2110 19584 2178 19640
rect 2234 19584 2302 19640
rect 2358 19584 2382 19640
rect 1906 19516 2382 19584
rect 1906 19460 1930 19516
rect 1986 19460 2054 19516
rect 2110 19460 2178 19516
rect 2234 19460 2302 19516
rect 2358 19460 2382 19516
rect 1906 19400 2382 19460
rect 86588 19640 87064 19708
rect 86588 19584 86612 19640
rect 86668 19584 86736 19640
rect 86792 19584 86860 19640
rect 86916 19584 86984 19640
rect 87040 19584 87064 19640
rect 86588 19516 87064 19584
rect 86588 19460 86612 19516
rect 86668 19460 86736 19516
rect 86792 19460 86860 19516
rect 86916 19460 86984 19516
rect 87040 19460 87064 19516
rect 86588 19392 87064 19460
rect 86588 19336 86612 19392
rect 86668 19336 86736 19392
rect 86792 19336 86860 19392
rect 86916 19336 86984 19392
rect 87040 19336 87064 19392
rect 86588 19324 87064 19336
rect 1106 18864 1582 18876
rect 1106 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1582 18864
rect 1106 18740 1582 18808
rect 1106 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1582 18740
rect 1106 18616 1582 18684
rect 1106 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1582 18616
rect 1106 18492 1582 18560
rect 1106 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1582 18492
rect 1106 18424 1582 18436
rect 85788 18864 86264 18876
rect 85788 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86264 18864
rect 85788 18740 86264 18808
rect 85788 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86264 18740
rect 85788 18616 86264 18684
rect 85788 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86264 18616
rect 85788 18492 86264 18560
rect 85788 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86264 18492
rect 85788 18424 86264 18436
rect 86588 17964 87064 17976
rect 86588 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87064 17964
rect 1906 17840 2382 17900
rect 1906 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2382 17840
rect 1906 17716 2382 17784
rect 1906 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2382 17716
rect 1906 17600 2382 17660
rect 86588 17840 87064 17908
rect 86588 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87064 17840
rect 86588 17716 87064 17784
rect 86588 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87064 17716
rect 86588 17592 87064 17660
rect 86588 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87064 17592
rect 86588 17524 87064 17536
rect 1106 17064 1582 17076
rect 1106 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1582 17064
rect 1106 16940 1582 17008
rect 1106 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1582 16940
rect 1106 16816 1582 16884
rect 1106 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1582 16816
rect 1106 16692 1582 16760
rect 1106 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1582 16692
rect 1106 16624 1582 16636
rect 85788 17064 86264 17076
rect 85788 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86264 17064
rect 85788 16940 86264 17008
rect 85788 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86264 16940
rect 85788 16816 86264 16884
rect 85788 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86264 16816
rect 85788 16692 86264 16760
rect 85788 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86264 16692
rect 85788 16624 86264 16636
rect 86588 16164 87064 16176
rect 86588 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87064 16164
rect 1906 16040 2382 16100
rect 1906 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2382 16040
rect 1906 15916 2382 15984
rect 1906 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2382 15916
rect 1906 15800 2382 15860
rect 86588 16040 87064 16108
rect 86588 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87064 16040
rect 86588 15916 87064 15984
rect 86588 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87064 15916
rect 86588 15792 87064 15860
rect 86588 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87064 15792
rect 86588 15724 87064 15736
rect 1106 15264 1582 15276
rect 1106 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1582 15264
rect 1106 15140 1582 15208
rect 1106 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1582 15140
rect 1106 15016 1582 15084
rect 1106 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1582 15016
rect 1106 14892 1582 14960
rect 1106 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1582 14892
rect 1106 14824 1582 14836
rect 85788 15264 86264 15276
rect 85788 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86264 15264
rect 85788 15140 86264 15208
rect 85788 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86264 15140
rect 85788 15016 86264 15084
rect 85788 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86264 15016
rect 85788 14892 86264 14960
rect 85788 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86264 14892
rect 85788 14824 86264 14836
rect 86588 14364 87064 14376
rect 86588 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87064 14364
rect 1906 14240 2382 14300
rect 1906 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2382 14240
rect 1906 14116 2382 14184
rect 1906 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2382 14116
rect 1906 14000 2382 14060
rect 86588 14240 87064 14308
rect 86588 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87064 14240
rect 86588 14116 87064 14184
rect 86588 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87064 14116
rect 86588 13992 87064 14060
rect 86588 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87064 13992
rect 86588 13924 87064 13936
rect 1106 13464 1582 13476
rect 1106 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1582 13464
rect 1106 13340 1582 13408
rect 1106 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1582 13340
rect 1106 13216 1582 13284
rect 1106 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1582 13216
rect 1106 13092 1582 13160
rect 1106 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1582 13092
rect 1106 13024 1582 13036
rect 85788 13464 86264 13476
rect 85788 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86264 13464
rect 85788 13340 86264 13408
rect 85788 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86264 13340
rect 85788 13216 86264 13284
rect 85788 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86264 13216
rect 85788 13092 86264 13160
rect 85788 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86264 13092
rect 85788 13024 86264 13036
rect 86588 12564 87064 12576
rect 86588 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87064 12564
rect 1906 12440 2382 12500
rect 1906 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2382 12440
rect 1906 12316 2382 12384
rect 1906 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2382 12316
rect 1906 12200 2382 12260
rect 86588 12440 87064 12508
rect 86588 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87064 12440
rect 86588 12316 87064 12384
rect 86588 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87064 12316
rect 86588 12192 87064 12260
rect 86588 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87064 12192
rect 86588 12124 87064 12136
rect 1106 11664 1582 11676
rect 1106 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1582 11664
rect 1106 11540 1582 11608
rect 1106 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1582 11540
rect 1106 11416 1582 11484
rect 1106 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1582 11416
rect 1106 11292 1582 11360
rect 1106 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1582 11292
rect 1106 11224 1582 11236
rect 85788 11664 86264 11676
rect 85788 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86264 11664
rect 85788 11540 86264 11608
rect 85788 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86264 11540
rect 85788 11416 86264 11484
rect 85788 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86264 11416
rect 85788 11292 86264 11360
rect 85788 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86264 11292
rect 85788 11224 86264 11236
rect 86588 10764 87064 10776
rect 86588 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87064 10764
rect 1906 10640 2382 10700
rect 1906 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2382 10640
rect 1906 10516 2382 10584
rect 1906 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2382 10516
rect 1906 10400 2382 10460
rect 86588 10640 87064 10708
rect 86588 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87064 10640
rect 86588 10516 87064 10584
rect 86588 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87064 10516
rect 86588 10392 87064 10460
rect 86588 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87064 10392
rect 86588 10324 87064 10336
rect 1106 9864 1582 9876
rect 1106 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1582 9864
rect 1106 9740 1582 9808
rect 1106 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1582 9740
rect 1106 9616 1582 9684
rect 1106 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1582 9616
rect 1106 9492 1582 9560
rect 1106 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1582 9492
rect 1106 9424 1582 9436
rect 85788 9864 86264 9876
rect 85788 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86264 9864
rect 85788 9740 86264 9808
rect 85788 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86264 9740
rect 85788 9616 86264 9684
rect 85788 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86264 9616
rect 85788 9492 86264 9560
rect 85788 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86264 9492
rect 85788 9424 86264 9436
rect 86588 8964 87064 8976
rect 86588 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87064 8964
rect 1906 8840 2382 8900
rect 1906 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2382 8840
rect 1906 8716 2382 8784
rect 1906 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2382 8716
rect 1906 8600 2382 8660
rect 86588 8840 87064 8908
rect 86588 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87064 8840
rect 86588 8716 87064 8784
rect 86588 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87064 8716
rect 86588 8592 87064 8660
rect 86588 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87064 8592
rect 86588 8524 87064 8536
rect 1106 8064 1582 8076
rect 1106 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1582 8064
rect 1106 7940 1582 8008
rect 1106 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1582 7940
rect 1106 7816 1582 7884
rect 1106 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1582 7816
rect 1106 7692 1582 7760
rect 1106 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1582 7692
rect 1106 7624 1582 7636
rect 85788 8064 86264 8076
rect 85788 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86264 8064
rect 85788 7940 86264 8008
rect 85788 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86264 7940
rect 85788 7816 86264 7884
rect 85788 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86264 7816
rect 85788 7692 86264 7760
rect 85788 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86264 7692
rect 85788 7624 86264 7636
rect 86588 7164 87064 7176
rect 86588 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87064 7164
rect 1906 7040 2382 7100
rect 1906 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2382 7040
rect 1906 6916 2382 6984
rect 1906 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2382 6916
rect 1906 6800 2382 6860
rect 86588 7040 87064 7108
rect 86588 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87064 7040
rect 86588 6916 87064 6984
rect 86588 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87064 6916
rect 86588 6792 87064 6860
rect 86588 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87064 6792
rect 86588 6724 87064 6736
rect 1106 6264 1582 6276
rect 1106 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1582 6264
rect 1106 6140 1582 6208
rect 1106 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1582 6140
rect 1106 6016 1582 6084
rect 1106 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1582 6016
rect 1106 5892 1582 5960
rect 1106 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1582 5892
rect 1106 5824 1582 5836
rect 85788 6264 86264 6276
rect 85788 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86264 6264
rect 85788 6140 86264 6208
rect 85788 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86264 6140
rect 85788 6016 86264 6084
rect 85788 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86264 6016
rect 85788 5892 86264 5960
rect 85788 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86264 5892
rect 85788 5824 86264 5836
rect 86588 5364 87064 5376
rect 86588 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87064 5364
rect 1906 5240 2382 5300
rect 1906 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2382 5240
rect 1906 5116 2382 5184
rect 1906 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2382 5116
rect 1906 5000 2382 5060
rect 86588 5240 87064 5308
rect 86588 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87064 5240
rect 86588 5116 87064 5184
rect 86588 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87064 5116
rect 86588 4992 87064 5060
rect 86588 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87064 4992
rect 86588 4924 87064 4936
rect 1106 4464 1582 4476
rect 1106 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1582 4464
rect 1106 4340 1582 4408
rect 1106 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1582 4340
rect 1106 4216 1582 4284
rect 1106 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1582 4216
rect 1106 4092 1582 4160
rect 1106 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1582 4092
rect 1106 4024 1582 4036
rect 85788 4464 86264 4476
rect 85788 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86264 4464
rect 85788 4340 86264 4408
rect 85788 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86264 4340
rect 85788 4216 86264 4284
rect 85788 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86264 4216
rect 85788 4092 86264 4160
rect 85788 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86264 4092
rect 85788 4024 86264 4036
rect 86588 3632 87064 3700
rect 86588 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87064 3632
rect 86588 3508 87064 3576
rect 1906 3440 2382 3500
rect 1906 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2382 3440
rect 1906 3316 2382 3384
rect 1906 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2382 3316
rect 1906 3200 2382 3260
rect 86588 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87064 3508
rect 86588 3384 87064 3452
rect 86588 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87064 3384
rect 86588 3260 87064 3328
rect 86588 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87064 3260
rect 86588 3136 87064 3204
<< via3 >>
rect 1901 95369 1957 95425
rect 1901 95245 1957 95301
rect 1901 95121 1957 95177
rect 1901 94997 1957 95053
rect 1901 94873 1957 94929
rect 1901 94749 1957 94805
rect 1901 94625 1957 94681
rect 1901 94501 1957 94557
rect 1901 94377 1957 94433
rect 1901 94253 1957 94309
rect 86550 95369 86606 95425
rect 86550 95245 86606 95301
rect 86550 95121 86606 95177
rect 86550 94997 86606 95053
rect 86550 94873 86606 94929
rect 86550 94749 86606 94805
rect 86550 94625 86606 94681
rect 86550 94501 86606 94557
rect 86550 94377 86606 94433
rect 86550 94253 86606 94309
rect 86674 95369 86730 95425
rect 86798 95369 86854 95425
rect 86922 95369 86978 95425
rect 87046 95369 87102 95425
rect 86674 95245 86730 95301
rect 86798 95245 86854 95301
rect 86922 95245 86978 95301
rect 87046 95245 87102 95301
rect 86674 95121 86730 95177
rect 86798 95121 86854 95177
rect 86922 95121 86978 95177
rect 87046 95121 87102 95177
rect 86674 94997 86730 95053
rect 86798 94997 86854 95053
rect 86922 94997 86978 95053
rect 87046 94997 87102 95053
rect 86674 94873 86730 94929
rect 86798 94873 86854 94929
rect 86922 94873 86978 94929
rect 87046 94873 87102 94929
rect 86674 94749 86730 94805
rect 86798 94749 86854 94805
rect 86922 94749 86978 94805
rect 87046 94749 87102 94805
rect 86674 94625 86730 94681
rect 86798 94625 86854 94681
rect 86922 94625 86978 94681
rect 87046 94625 87102 94681
rect 86674 94501 86730 94557
rect 86798 94501 86854 94557
rect 86922 94501 86978 94557
rect 87046 94501 87102 94557
rect 86674 94377 86730 94433
rect 86798 94377 86854 94433
rect 86922 94377 86978 94433
rect 87046 94377 87102 94433
rect 86674 94253 86730 94309
rect 86798 94253 86854 94309
rect 86922 94253 86978 94309
rect 87046 94253 87102 94309
rect 86550 92135 86606 92191
rect 86550 92011 86606 92067
rect 86550 91887 86606 91943
rect 86550 91763 86606 91819
rect 86674 92135 86730 92191
rect 86798 92135 86854 92191
rect 86922 92135 86978 92191
rect 87046 92135 87102 92191
rect 86674 92011 86730 92067
rect 86798 92011 86854 92067
rect 86922 92011 86978 92067
rect 87046 92011 87102 92067
rect 86674 91887 86730 91943
rect 86798 91887 86854 91943
rect 86922 91887 86978 91943
rect 87046 91887 87102 91943
rect 86674 91763 86730 91819
rect 86798 91763 86854 91819
rect 86922 91763 86978 91819
rect 87046 91763 87102 91819
rect 86550 91639 86606 91695
rect 86550 91515 86606 91571
rect 86550 91391 86606 91447
rect 86550 91267 86606 91323
rect 86674 91639 86730 91695
rect 86798 91639 86854 91695
rect 86922 91639 86978 91695
rect 87046 91639 87102 91695
rect 86674 91515 86730 91571
rect 86798 91515 86854 91571
rect 86922 91515 86978 91571
rect 87046 91515 87102 91571
rect 86674 91391 86730 91447
rect 86798 91391 86854 91447
rect 86922 91391 86978 91447
rect 87046 91391 87102 91447
rect 86674 91267 86730 91323
rect 86798 91267 86854 91323
rect 86922 91267 86978 91323
rect 87046 91267 87102 91323
rect 86550 91143 86606 91199
rect 86550 91019 86606 91075
rect 1930 90845 1986 90901
rect 2054 90845 2110 90901
rect 2178 90845 2234 90901
rect 2302 90845 2358 90901
rect 1930 90721 1986 90777
rect 2054 90721 2110 90777
rect 2178 90721 2234 90777
rect 2302 90721 2358 90777
rect 86550 90895 86606 90951
rect 86550 90771 86606 90827
rect 86674 91143 86730 91199
rect 86798 91143 86854 91199
rect 86922 91143 86978 91199
rect 87046 91143 87102 91199
rect 86674 91019 86730 91075
rect 86798 91019 86854 91075
rect 86922 91019 86978 91075
rect 87046 91019 87102 91075
rect 86674 90895 86730 90951
rect 86798 90895 86854 90951
rect 86922 90895 86978 90951
rect 87046 90895 87102 90951
rect 86674 90771 86730 90827
rect 86798 90771 86854 90827
rect 86922 90771 86978 90827
rect 87046 90771 87102 90827
rect 1930 90597 1986 90653
rect 2054 90597 2110 90653
rect 2178 90597 2234 90653
rect 2302 90597 2358 90653
rect 1930 90473 1986 90529
rect 2054 90473 2110 90529
rect 2178 90473 2234 90529
rect 2302 90473 2358 90529
rect 86550 90647 86606 90703
rect 86550 90523 86606 90579
rect 86550 90399 86606 90455
rect 86674 90647 86730 90703
rect 86798 90647 86854 90703
rect 86922 90647 86978 90703
rect 87046 90647 87102 90703
rect 86674 90523 86730 90579
rect 86798 90523 86854 90579
rect 86922 90523 86978 90579
rect 87046 90523 87102 90579
rect 86674 90399 86730 90455
rect 86798 90399 86854 90455
rect 86922 90399 86978 90455
rect 87046 90399 87102 90455
rect 85750 89735 85806 89791
rect 85750 89611 85806 89667
rect 85750 89487 85806 89543
rect 85750 89363 85806 89419
rect 85874 89735 85930 89791
rect 85998 89735 86054 89791
rect 86122 89735 86178 89791
rect 86246 89735 86302 89791
rect 85874 89611 85930 89667
rect 85998 89611 86054 89667
rect 86122 89611 86178 89667
rect 86246 89611 86302 89667
rect 85874 89487 85930 89543
rect 85998 89487 86054 89543
rect 86122 89487 86178 89543
rect 86246 89487 86302 89543
rect 85874 89363 85930 89419
rect 85998 89363 86054 89419
rect 86122 89363 86178 89419
rect 86246 89363 86302 89419
rect 85750 89239 85806 89295
rect 85750 89115 85806 89171
rect 85750 88991 85806 89047
rect 85750 88867 85806 88923
rect 85874 89239 85930 89295
rect 85998 89239 86054 89295
rect 86122 89239 86178 89295
rect 86246 89239 86302 89295
rect 85874 89115 85930 89171
rect 85998 89115 86054 89171
rect 86122 89115 86178 89171
rect 86246 89115 86302 89171
rect 85874 88991 85930 89047
rect 85998 88991 86054 89047
rect 86122 88991 86178 89047
rect 86246 88991 86302 89047
rect 85874 88867 85930 88923
rect 85998 88867 86054 88923
rect 86122 88867 86178 88923
rect 86246 88867 86302 88923
rect 85750 88743 85806 88799
rect 85750 88619 85806 88675
rect 85750 88495 85806 88551
rect 85874 88743 85930 88799
rect 85998 88743 86054 88799
rect 86122 88743 86178 88799
rect 86246 88743 86302 88799
rect 85874 88619 85930 88675
rect 85998 88619 86054 88675
rect 86122 88619 86178 88675
rect 86246 88619 86302 88675
rect 85874 88495 85930 88551
rect 85998 88495 86054 88551
rect 86122 88495 86178 88551
rect 86246 88495 86302 88551
rect 1068 85833 1124 85889
rect 1068 85709 1124 85765
rect 1068 85585 1124 85641
rect 1068 85461 1124 85517
rect 1068 85337 1124 85393
rect 1068 85213 1124 85269
rect 1068 85089 1124 85145
rect 1068 84965 1124 85021
rect 1068 84841 1124 84897
rect 1068 84717 1124 84773
rect 1068 84593 1124 84649
rect 1068 84469 1124 84525
rect 1068 84345 1124 84401
rect 1068 84221 1124 84277
rect 1068 84097 1124 84153
rect 1068 83973 1124 84029
rect 1068 83849 1124 83905
rect 1192 85833 1248 85889
rect 1316 85833 1372 85889
rect 1440 85833 1496 85889
rect 1564 85833 1620 85889
rect 1192 85709 1248 85765
rect 1316 85709 1372 85765
rect 1440 85709 1496 85765
rect 1564 85709 1620 85765
rect 1192 85585 1248 85641
rect 1316 85585 1372 85641
rect 1440 85585 1496 85641
rect 1564 85585 1620 85641
rect 1192 85461 1248 85517
rect 1316 85461 1372 85517
rect 1440 85461 1496 85517
rect 1564 85461 1620 85517
rect 1192 85337 1248 85393
rect 1316 85337 1372 85393
rect 1440 85337 1496 85393
rect 1564 85337 1620 85393
rect 1192 85213 1248 85269
rect 1316 85213 1372 85269
rect 1440 85213 1496 85269
rect 1564 85213 1620 85269
rect 1192 85089 1248 85145
rect 1316 85089 1372 85145
rect 1440 85089 1496 85145
rect 1564 85089 1620 85145
rect 1192 84965 1248 85021
rect 1316 84965 1372 85021
rect 1440 84965 1496 85021
rect 1564 84965 1620 85021
rect 1192 84841 1248 84897
rect 1316 84841 1372 84897
rect 1440 84841 1496 84897
rect 1564 84841 1620 84897
rect 1192 84717 1248 84773
rect 1316 84717 1372 84773
rect 1440 84717 1496 84773
rect 1564 84717 1620 84773
rect 1192 84593 1248 84649
rect 1316 84593 1372 84649
rect 1440 84593 1496 84649
rect 1564 84593 1620 84649
rect 1192 84469 1248 84525
rect 1316 84469 1372 84525
rect 1440 84469 1496 84525
rect 1564 84469 1620 84525
rect 1192 84345 1248 84401
rect 1316 84345 1372 84401
rect 1440 84345 1496 84401
rect 1564 84345 1620 84401
rect 1192 84221 1248 84277
rect 1316 84221 1372 84277
rect 1440 84221 1496 84277
rect 1564 84221 1620 84277
rect 1192 84097 1248 84153
rect 1316 84097 1372 84153
rect 1440 84097 1496 84153
rect 1564 84097 1620 84153
rect 1192 83973 1248 84029
rect 1316 83973 1372 84029
rect 1440 83973 1496 84029
rect 1564 83973 1620 84029
rect 1192 83849 1248 83905
rect 1316 83849 1372 83905
rect 1440 83849 1496 83905
rect 1564 83849 1620 83905
rect 85750 85833 85806 85889
rect 85750 85709 85806 85765
rect 85750 85585 85806 85641
rect 85750 85461 85806 85517
rect 85750 85337 85806 85393
rect 85750 85213 85806 85269
rect 85750 85089 85806 85145
rect 85750 84965 85806 85021
rect 85750 84841 85806 84897
rect 85750 84717 85806 84773
rect 85750 84593 85806 84649
rect 85750 84469 85806 84525
rect 85750 84345 85806 84401
rect 85750 84221 85806 84277
rect 85750 84097 85806 84153
rect 85750 83973 85806 84029
rect 85750 83849 85806 83905
rect 85874 85833 85930 85889
rect 85998 85833 86054 85889
rect 86122 85833 86178 85889
rect 86246 85833 86302 85889
rect 85874 85709 85930 85765
rect 85998 85709 86054 85765
rect 86122 85709 86178 85765
rect 86246 85709 86302 85765
rect 85874 85585 85930 85641
rect 85998 85585 86054 85641
rect 86122 85585 86178 85641
rect 86246 85585 86302 85641
rect 85874 85461 85930 85517
rect 85998 85461 86054 85517
rect 86122 85461 86178 85517
rect 86246 85461 86302 85517
rect 85874 85337 85930 85393
rect 85998 85337 86054 85393
rect 86122 85337 86178 85393
rect 86246 85337 86302 85393
rect 85874 85213 85930 85269
rect 85998 85213 86054 85269
rect 86122 85213 86178 85269
rect 86246 85213 86302 85269
rect 85874 85089 85930 85145
rect 85998 85089 86054 85145
rect 86122 85089 86178 85145
rect 86246 85089 86302 85145
rect 85874 84965 85930 85021
rect 85998 84965 86054 85021
rect 86122 84965 86178 85021
rect 86246 84965 86302 85021
rect 85874 84841 85930 84897
rect 85998 84841 86054 84897
rect 86122 84841 86178 84897
rect 86246 84841 86302 84897
rect 85874 84717 85930 84773
rect 85998 84717 86054 84773
rect 86122 84717 86178 84773
rect 86246 84717 86302 84773
rect 85874 84593 85930 84649
rect 85998 84593 86054 84649
rect 86122 84593 86178 84649
rect 86246 84593 86302 84649
rect 85874 84469 85930 84525
rect 85998 84469 86054 84525
rect 86122 84469 86178 84525
rect 86246 84469 86302 84525
rect 85874 84345 85930 84401
rect 85998 84345 86054 84401
rect 86122 84345 86178 84401
rect 86246 84345 86302 84401
rect 85874 84221 85930 84277
rect 85998 84221 86054 84277
rect 86122 84221 86178 84277
rect 86246 84221 86302 84277
rect 85874 84097 85930 84153
rect 85998 84097 86054 84153
rect 86122 84097 86178 84153
rect 86246 84097 86302 84153
rect 85874 83973 85930 84029
rect 85998 83973 86054 84029
rect 86122 83973 86178 84029
rect 86246 83973 86302 84029
rect 85874 83849 85930 83905
rect 85998 83849 86054 83905
rect 86122 83849 86178 83905
rect 86246 83849 86302 83905
rect 1868 83531 1924 83587
rect 1868 83407 1924 83463
rect 1868 83283 1924 83339
rect 1868 83159 1924 83215
rect 1868 83035 1924 83091
rect 1868 82911 1924 82967
rect 1868 82787 1924 82843
rect 1868 82663 1924 82719
rect 1868 82539 1924 82595
rect 1868 82415 1924 82471
rect 1868 82291 1924 82347
rect 1868 82167 1924 82223
rect 1868 82043 1924 82099
rect 1868 81919 1924 81975
rect 1868 81795 1924 81851
rect 1868 81671 1924 81727
rect 1868 81547 1924 81603
rect 1868 81423 1924 81479
rect 1868 81299 1924 81355
rect 1868 81175 1924 81231
rect 1868 81051 1924 81107
rect 1868 80927 1924 80983
rect 1868 80803 1924 80859
rect 1868 80679 1924 80735
rect 1868 80555 1924 80611
rect 1868 80431 1924 80487
rect 1868 80307 1924 80363
rect 1992 83531 2048 83587
rect 2116 83531 2172 83587
rect 2240 83531 2296 83587
rect 2364 83531 2420 83587
rect 1992 83407 2048 83463
rect 2116 83407 2172 83463
rect 2240 83407 2296 83463
rect 2364 83407 2420 83463
rect 1992 83283 2048 83339
rect 2116 83283 2172 83339
rect 2240 83283 2296 83339
rect 2364 83283 2420 83339
rect 1992 83159 2048 83215
rect 2116 83159 2172 83215
rect 2240 83159 2296 83215
rect 2364 83159 2420 83215
rect 1992 83035 2048 83091
rect 2116 83035 2172 83091
rect 2240 83035 2296 83091
rect 2364 83035 2420 83091
rect 1992 82911 2048 82967
rect 2116 82911 2172 82967
rect 2240 82911 2296 82967
rect 2364 82911 2420 82967
rect 1992 82787 2048 82843
rect 2116 82787 2172 82843
rect 2240 82787 2296 82843
rect 2364 82787 2420 82843
rect 1992 82663 2048 82719
rect 2116 82663 2172 82719
rect 2240 82663 2296 82719
rect 2364 82663 2420 82719
rect 1992 82539 2048 82595
rect 2116 82539 2172 82595
rect 2240 82539 2296 82595
rect 2364 82539 2420 82595
rect 1992 82415 2048 82471
rect 2116 82415 2172 82471
rect 2240 82415 2296 82471
rect 2364 82415 2420 82471
rect 1992 82291 2048 82347
rect 2116 82291 2172 82347
rect 2240 82291 2296 82347
rect 2364 82291 2420 82347
rect 1992 82167 2048 82223
rect 2116 82167 2172 82223
rect 2240 82167 2296 82223
rect 2364 82167 2420 82223
rect 1992 82043 2048 82099
rect 2116 82043 2172 82099
rect 2240 82043 2296 82099
rect 2364 82043 2420 82099
rect 1992 81919 2048 81975
rect 2116 81919 2172 81975
rect 2240 81919 2296 81975
rect 2364 81919 2420 81975
rect 1992 81795 2048 81851
rect 2116 81795 2172 81851
rect 2240 81795 2296 81851
rect 2364 81795 2420 81851
rect 1992 81671 2048 81727
rect 2116 81671 2172 81727
rect 2240 81671 2296 81727
rect 2364 81671 2420 81727
rect 1992 81547 2048 81603
rect 2116 81547 2172 81603
rect 2240 81547 2296 81603
rect 2364 81547 2420 81603
rect 1992 81423 2048 81479
rect 2116 81423 2172 81479
rect 2240 81423 2296 81479
rect 2364 81423 2420 81479
rect 1992 81299 2048 81355
rect 2116 81299 2172 81355
rect 2240 81299 2296 81355
rect 2364 81299 2420 81355
rect 1992 81175 2048 81231
rect 2116 81175 2172 81231
rect 2240 81175 2296 81231
rect 2364 81175 2420 81231
rect 1992 81051 2048 81107
rect 2116 81051 2172 81107
rect 2240 81051 2296 81107
rect 2364 81051 2420 81107
rect 1992 80927 2048 80983
rect 2116 80927 2172 80983
rect 2240 80927 2296 80983
rect 2364 80927 2420 80983
rect 1992 80803 2048 80859
rect 2116 80803 2172 80859
rect 2240 80803 2296 80859
rect 2364 80803 2420 80859
rect 1992 80679 2048 80735
rect 2116 80679 2172 80735
rect 2240 80679 2296 80735
rect 2364 80679 2420 80735
rect 1992 80555 2048 80611
rect 2116 80555 2172 80611
rect 2240 80555 2296 80611
rect 2364 80555 2420 80611
rect 1992 80431 2048 80487
rect 2116 80431 2172 80487
rect 2240 80431 2296 80487
rect 2364 80431 2420 80487
rect 1992 80307 2048 80363
rect 2116 80307 2172 80363
rect 2240 80307 2296 80363
rect 2364 80307 2420 80363
rect 86550 83531 86606 83587
rect 86550 83407 86606 83463
rect 86550 83283 86606 83339
rect 86550 83159 86606 83215
rect 86550 83035 86606 83091
rect 86550 82911 86606 82967
rect 86550 82787 86606 82843
rect 86550 82663 86606 82719
rect 86550 82539 86606 82595
rect 86550 82415 86606 82471
rect 86550 82291 86606 82347
rect 86550 82167 86606 82223
rect 86550 82043 86606 82099
rect 86550 81919 86606 81975
rect 86550 81795 86606 81851
rect 86550 81671 86606 81727
rect 86550 81547 86606 81603
rect 86550 81423 86606 81479
rect 86550 81299 86606 81355
rect 86550 81175 86606 81231
rect 86550 81051 86606 81107
rect 86550 80927 86606 80983
rect 86550 80803 86606 80859
rect 86550 80679 86606 80735
rect 86550 80555 86606 80611
rect 86550 80431 86606 80487
rect 86550 80307 86606 80363
rect 86674 83531 86730 83587
rect 86798 83531 86854 83587
rect 86922 83531 86978 83587
rect 87046 83531 87102 83587
rect 86674 83407 86730 83463
rect 86798 83407 86854 83463
rect 86922 83407 86978 83463
rect 87046 83407 87102 83463
rect 86674 83283 86730 83339
rect 86798 83283 86854 83339
rect 86922 83283 86978 83339
rect 87046 83283 87102 83339
rect 86674 83159 86730 83215
rect 86798 83159 86854 83215
rect 86922 83159 86978 83215
rect 87046 83159 87102 83215
rect 86674 83035 86730 83091
rect 86798 83035 86854 83091
rect 86922 83035 86978 83091
rect 87046 83035 87102 83091
rect 86674 82911 86730 82967
rect 86798 82911 86854 82967
rect 86922 82911 86978 82967
rect 87046 82911 87102 82967
rect 86674 82787 86730 82843
rect 86798 82787 86854 82843
rect 86922 82787 86978 82843
rect 87046 82787 87102 82843
rect 86674 82663 86730 82719
rect 86798 82663 86854 82719
rect 86922 82663 86978 82719
rect 87046 82663 87102 82719
rect 86674 82539 86730 82595
rect 86798 82539 86854 82595
rect 86922 82539 86978 82595
rect 87046 82539 87102 82595
rect 86674 82415 86730 82471
rect 86798 82415 86854 82471
rect 86922 82415 86978 82471
rect 87046 82415 87102 82471
rect 86674 82291 86730 82347
rect 86798 82291 86854 82347
rect 86922 82291 86978 82347
rect 87046 82291 87102 82347
rect 86674 82167 86730 82223
rect 86798 82167 86854 82223
rect 86922 82167 86978 82223
rect 87046 82167 87102 82223
rect 86674 82043 86730 82099
rect 86798 82043 86854 82099
rect 86922 82043 86978 82099
rect 87046 82043 87102 82099
rect 86674 81919 86730 81975
rect 86798 81919 86854 81975
rect 86922 81919 86978 81975
rect 87046 81919 87102 81975
rect 86674 81795 86730 81851
rect 86798 81795 86854 81851
rect 86922 81795 86978 81851
rect 87046 81795 87102 81851
rect 86674 81671 86730 81727
rect 86798 81671 86854 81727
rect 86922 81671 86978 81727
rect 87046 81671 87102 81727
rect 86674 81547 86730 81603
rect 86798 81547 86854 81603
rect 86922 81547 86978 81603
rect 87046 81547 87102 81603
rect 86674 81423 86730 81479
rect 86798 81423 86854 81479
rect 86922 81423 86978 81479
rect 87046 81423 87102 81479
rect 86674 81299 86730 81355
rect 86798 81299 86854 81355
rect 86922 81299 86978 81355
rect 87046 81299 87102 81355
rect 86674 81175 86730 81231
rect 86798 81175 86854 81231
rect 86922 81175 86978 81231
rect 87046 81175 87102 81231
rect 86674 81051 86730 81107
rect 86798 81051 86854 81107
rect 86922 81051 86978 81107
rect 87046 81051 87102 81107
rect 86674 80927 86730 80983
rect 86798 80927 86854 80983
rect 86922 80927 86978 80983
rect 87046 80927 87102 80983
rect 86674 80803 86730 80859
rect 86798 80803 86854 80859
rect 86922 80803 86978 80859
rect 87046 80803 87102 80859
rect 86674 80679 86730 80735
rect 86798 80679 86854 80735
rect 86922 80679 86978 80735
rect 87046 80679 87102 80735
rect 86674 80555 86730 80611
rect 86798 80555 86854 80611
rect 86922 80555 86978 80611
rect 87046 80555 87102 80611
rect 86674 80431 86730 80487
rect 86798 80431 86854 80487
rect 86922 80431 86978 80487
rect 87046 80431 87102 80487
rect 86674 80307 86730 80363
rect 86798 80307 86854 80363
rect 86922 80307 86978 80363
rect 87046 80307 87102 80363
rect 86550 76600 86606 76656
rect 86550 76476 86606 76532
rect 86550 76352 86606 76408
rect 86550 76228 86606 76284
rect 86550 76104 86606 76160
rect 86550 75980 86606 76036
rect 86550 75856 86606 75912
rect 86550 75732 86606 75788
rect 86674 76600 86730 76656
rect 86798 76600 86854 76656
rect 86922 76600 86978 76656
rect 87046 76600 87102 76656
rect 86674 76476 86730 76532
rect 86798 76476 86854 76532
rect 86922 76476 86978 76532
rect 87046 76476 87102 76532
rect 86674 76352 86730 76408
rect 86798 76352 86854 76408
rect 86922 76352 86978 76408
rect 87046 76352 87102 76408
rect 86674 76228 86730 76284
rect 86798 76228 86854 76284
rect 86922 76228 86978 76284
rect 87046 76228 87102 76284
rect 86674 76104 86730 76160
rect 86798 76104 86854 76160
rect 86922 76104 86978 76160
rect 87046 76104 87102 76160
rect 86674 75980 86730 76036
rect 86798 75980 86854 76036
rect 86922 75980 86978 76036
rect 87046 75980 87102 76036
rect 86674 75856 86730 75912
rect 86798 75856 86854 75912
rect 86922 75856 86978 75912
rect 87046 75856 87102 75912
rect 86674 75732 86730 75788
rect 86798 75732 86854 75788
rect 86922 75732 86978 75788
rect 87046 75732 87102 75788
rect 1068 74944 1124 75000
rect 1068 74820 1124 74876
rect 1068 74696 1124 74752
rect 1068 74572 1124 74628
rect 1068 74448 1124 74504
rect 1068 74324 1124 74380
rect 1068 74200 1124 74256
rect 1068 74076 1124 74132
rect 1192 74944 1248 75000
rect 1316 74944 1372 75000
rect 1440 74944 1496 75000
rect 1564 74944 1620 75000
rect 1192 74820 1248 74876
rect 1316 74820 1372 74876
rect 1440 74820 1496 74876
rect 1564 74820 1620 74876
rect 1192 74696 1248 74752
rect 1316 74696 1372 74752
rect 1440 74696 1496 74752
rect 1564 74696 1620 74752
rect 1192 74572 1248 74628
rect 1316 74572 1372 74628
rect 1440 74572 1496 74628
rect 1564 74572 1620 74628
rect 1192 74448 1248 74504
rect 1316 74448 1372 74504
rect 1440 74448 1496 74504
rect 1564 74448 1620 74504
rect 1192 74324 1248 74380
rect 1316 74324 1372 74380
rect 1440 74324 1496 74380
rect 1564 74324 1620 74380
rect 1192 74200 1248 74256
rect 1316 74200 1372 74256
rect 1440 74200 1496 74256
rect 1564 74200 1620 74256
rect 1192 74076 1248 74132
rect 1316 74076 1372 74132
rect 1440 74076 1496 74132
rect 1564 74076 1620 74132
rect 85750 74944 85806 75000
rect 85750 74820 85806 74876
rect 85750 74696 85806 74752
rect 85750 74572 85806 74628
rect 85750 74448 85806 74504
rect 85750 74324 85806 74380
rect 85750 74200 85806 74256
rect 85750 74076 85806 74132
rect 85874 74944 85930 75000
rect 85998 74944 86054 75000
rect 86122 74944 86178 75000
rect 86246 74944 86302 75000
rect 85874 74820 85930 74876
rect 85998 74820 86054 74876
rect 86122 74820 86178 74876
rect 86246 74820 86302 74876
rect 85874 74696 85930 74752
rect 85998 74696 86054 74752
rect 86122 74696 86178 74752
rect 86246 74696 86302 74752
rect 85874 74572 85930 74628
rect 85998 74572 86054 74628
rect 86122 74572 86178 74628
rect 86246 74572 86302 74628
rect 85874 74448 85930 74504
rect 85998 74448 86054 74504
rect 86122 74448 86178 74504
rect 86246 74448 86302 74504
rect 85874 74324 85930 74380
rect 85998 74324 86054 74380
rect 86122 74324 86178 74380
rect 86246 74324 86302 74380
rect 85874 74200 85930 74256
rect 85998 74200 86054 74256
rect 86122 74200 86178 74256
rect 86246 74200 86302 74256
rect 85874 74076 85930 74132
rect 85998 74076 86054 74132
rect 86122 74076 86178 74132
rect 86246 74076 86302 74132
rect 1930 63358 1986 63414
rect 2054 63358 2110 63414
rect 2178 63358 2234 63414
rect 2302 63358 2358 63414
rect 1930 63234 1986 63290
rect 2054 63234 2110 63290
rect 2178 63234 2234 63290
rect 2302 63234 2358 63290
rect 1930 63110 1986 63166
rect 2054 63110 2110 63166
rect 2178 63110 2234 63166
rect 2302 63110 2358 63166
rect 1930 62986 1986 63042
rect 2054 62986 2110 63042
rect 2178 62986 2234 63042
rect 2302 62986 2358 63042
rect 86612 63203 86668 63259
rect 86736 63203 86792 63259
rect 86860 63203 86916 63259
rect 86984 63203 87040 63259
rect 86612 63079 86668 63135
rect 86736 63079 86792 63135
rect 86860 63079 86916 63135
rect 86984 63079 87040 63135
rect 86612 62955 86668 63011
rect 86736 62955 86792 63011
rect 86860 62955 86916 63011
rect 86984 62955 87040 63011
rect 1930 62784 1986 62840
rect 2054 62784 2110 62840
rect 2178 62784 2234 62840
rect 2302 62784 2358 62840
rect 86612 62831 86668 62887
rect 86736 62831 86792 62887
rect 86860 62831 86916 62887
rect 86984 62831 87040 62887
rect 1930 62660 1986 62716
rect 2054 62660 2110 62716
rect 2178 62660 2234 62716
rect 2302 62660 2358 62716
rect 1130 62008 1186 62064
rect 1254 62008 1310 62064
rect 1378 62008 1434 62064
rect 1502 62008 1558 62064
rect 1130 61884 1186 61940
rect 1254 61884 1310 61940
rect 1378 61884 1434 61940
rect 1502 61884 1558 61940
rect 1130 61760 1186 61816
rect 1254 61760 1310 61816
rect 1378 61760 1434 61816
rect 1502 61760 1558 61816
rect 1130 61636 1186 61692
rect 1254 61636 1310 61692
rect 1378 61636 1434 61692
rect 1502 61636 1558 61692
rect 85812 62008 85868 62064
rect 85936 62008 85992 62064
rect 86060 62008 86116 62064
rect 86184 62008 86240 62064
rect 85812 61884 85868 61940
rect 85936 61884 85992 61940
rect 86060 61884 86116 61940
rect 86184 61884 86240 61940
rect 85812 61760 85868 61816
rect 85936 61760 85992 61816
rect 86060 61760 86116 61816
rect 86184 61760 86240 61816
rect 85812 61636 85868 61692
rect 85936 61636 85992 61692
rect 86060 61636 86116 61692
rect 86184 61636 86240 61692
rect 86612 61108 86668 61164
rect 86736 61108 86792 61164
rect 86860 61108 86916 61164
rect 86984 61108 87040 61164
rect 1930 60984 1986 61040
rect 2054 60984 2110 61040
rect 2178 60984 2234 61040
rect 2302 60984 2358 61040
rect 1930 60860 1986 60916
rect 2054 60860 2110 60916
rect 2178 60860 2234 60916
rect 2302 60860 2358 60916
rect 86612 60984 86668 61040
rect 86736 60984 86792 61040
rect 86860 60984 86916 61040
rect 86984 60984 87040 61040
rect 86612 60860 86668 60916
rect 86736 60860 86792 60916
rect 86860 60860 86916 60916
rect 86984 60860 87040 60916
rect 86612 60736 86668 60792
rect 86736 60736 86792 60792
rect 86860 60736 86916 60792
rect 86984 60736 87040 60792
rect 1130 60208 1186 60264
rect 1254 60208 1310 60264
rect 1378 60208 1434 60264
rect 1502 60208 1558 60264
rect 1130 60084 1186 60140
rect 1254 60084 1310 60140
rect 1378 60084 1434 60140
rect 1502 60084 1558 60140
rect 1130 59960 1186 60016
rect 1254 59960 1310 60016
rect 1378 59960 1434 60016
rect 1502 59960 1558 60016
rect 1130 59836 1186 59892
rect 1254 59836 1310 59892
rect 1378 59836 1434 59892
rect 1502 59836 1558 59892
rect 85812 60208 85868 60264
rect 85936 60208 85992 60264
rect 86060 60208 86116 60264
rect 86184 60208 86240 60264
rect 85812 60084 85868 60140
rect 85936 60084 85992 60140
rect 86060 60084 86116 60140
rect 86184 60084 86240 60140
rect 85812 59960 85868 60016
rect 85936 59960 85992 60016
rect 86060 59960 86116 60016
rect 86184 59960 86240 60016
rect 85812 59836 85868 59892
rect 85936 59836 85992 59892
rect 86060 59836 86116 59892
rect 86184 59836 86240 59892
rect 86612 59308 86668 59364
rect 86736 59308 86792 59364
rect 86860 59308 86916 59364
rect 86984 59308 87040 59364
rect 1930 59184 1986 59240
rect 2054 59184 2110 59240
rect 2178 59184 2234 59240
rect 2302 59184 2358 59240
rect 1930 59060 1986 59116
rect 2054 59060 2110 59116
rect 2178 59060 2234 59116
rect 2302 59060 2358 59116
rect 86612 59184 86668 59240
rect 86736 59184 86792 59240
rect 86860 59184 86916 59240
rect 86984 59184 87040 59240
rect 86612 59060 86668 59116
rect 86736 59060 86792 59116
rect 86860 59060 86916 59116
rect 86984 59060 87040 59116
rect 86612 58936 86668 58992
rect 86736 58936 86792 58992
rect 86860 58936 86916 58992
rect 86984 58936 87040 58992
rect 1130 58408 1186 58464
rect 1254 58408 1310 58464
rect 1378 58408 1434 58464
rect 1502 58408 1558 58464
rect 1130 58284 1186 58340
rect 1254 58284 1310 58340
rect 1378 58284 1434 58340
rect 1502 58284 1558 58340
rect 1130 58160 1186 58216
rect 1254 58160 1310 58216
rect 1378 58160 1434 58216
rect 1502 58160 1558 58216
rect 1130 58036 1186 58092
rect 1254 58036 1310 58092
rect 1378 58036 1434 58092
rect 1502 58036 1558 58092
rect 85812 58408 85868 58464
rect 85936 58408 85992 58464
rect 86060 58408 86116 58464
rect 86184 58408 86240 58464
rect 85812 58284 85868 58340
rect 85936 58284 85992 58340
rect 86060 58284 86116 58340
rect 86184 58284 86240 58340
rect 85812 58160 85868 58216
rect 85936 58160 85992 58216
rect 86060 58160 86116 58216
rect 86184 58160 86240 58216
rect 85812 58036 85868 58092
rect 85936 58036 85992 58092
rect 86060 58036 86116 58092
rect 86184 58036 86240 58092
rect 86612 57508 86668 57564
rect 86736 57508 86792 57564
rect 86860 57508 86916 57564
rect 86984 57508 87040 57564
rect 1930 57384 1986 57440
rect 2054 57384 2110 57440
rect 2178 57384 2234 57440
rect 2302 57384 2358 57440
rect 1930 57260 1986 57316
rect 2054 57260 2110 57316
rect 2178 57260 2234 57316
rect 2302 57260 2358 57316
rect 86612 57384 86668 57440
rect 86736 57384 86792 57440
rect 86860 57384 86916 57440
rect 86984 57384 87040 57440
rect 86612 57260 86668 57316
rect 86736 57260 86792 57316
rect 86860 57260 86916 57316
rect 86984 57260 87040 57316
rect 86612 57136 86668 57192
rect 86736 57136 86792 57192
rect 86860 57136 86916 57192
rect 86984 57136 87040 57192
rect 1130 56608 1186 56664
rect 1254 56608 1310 56664
rect 1378 56608 1434 56664
rect 1502 56608 1558 56664
rect 1130 56484 1186 56540
rect 1254 56484 1310 56540
rect 1378 56484 1434 56540
rect 1502 56484 1558 56540
rect 1130 56360 1186 56416
rect 1254 56360 1310 56416
rect 1378 56360 1434 56416
rect 1502 56360 1558 56416
rect 1130 56236 1186 56292
rect 1254 56236 1310 56292
rect 1378 56236 1434 56292
rect 1502 56236 1558 56292
rect 85812 56608 85868 56664
rect 85936 56608 85992 56664
rect 86060 56608 86116 56664
rect 86184 56608 86240 56664
rect 85812 56484 85868 56540
rect 85936 56484 85992 56540
rect 86060 56484 86116 56540
rect 86184 56484 86240 56540
rect 85812 56360 85868 56416
rect 85936 56360 85992 56416
rect 86060 56360 86116 56416
rect 86184 56360 86240 56416
rect 85812 56236 85868 56292
rect 85936 56236 85992 56292
rect 86060 56236 86116 56292
rect 86184 56236 86240 56292
rect 86612 55708 86668 55764
rect 86736 55708 86792 55764
rect 86860 55708 86916 55764
rect 86984 55708 87040 55764
rect 1930 55584 1986 55640
rect 2054 55584 2110 55640
rect 2178 55584 2234 55640
rect 2302 55584 2358 55640
rect 1930 55460 1986 55516
rect 2054 55460 2110 55516
rect 2178 55460 2234 55516
rect 2302 55460 2358 55516
rect 86612 55584 86668 55640
rect 86736 55584 86792 55640
rect 86860 55584 86916 55640
rect 86984 55584 87040 55640
rect 86612 55460 86668 55516
rect 86736 55460 86792 55516
rect 86860 55460 86916 55516
rect 86984 55460 87040 55516
rect 86612 55336 86668 55392
rect 86736 55336 86792 55392
rect 86860 55336 86916 55392
rect 86984 55336 87040 55392
rect 1130 54808 1186 54864
rect 1254 54808 1310 54864
rect 1378 54808 1434 54864
rect 1502 54808 1558 54864
rect 1130 54684 1186 54740
rect 1254 54684 1310 54740
rect 1378 54684 1434 54740
rect 1502 54684 1558 54740
rect 1130 54560 1186 54616
rect 1254 54560 1310 54616
rect 1378 54560 1434 54616
rect 1502 54560 1558 54616
rect 1130 54436 1186 54492
rect 1254 54436 1310 54492
rect 1378 54436 1434 54492
rect 1502 54436 1558 54492
rect 85812 54808 85868 54864
rect 85936 54808 85992 54864
rect 86060 54808 86116 54864
rect 86184 54808 86240 54864
rect 85812 54684 85868 54740
rect 85936 54684 85992 54740
rect 86060 54684 86116 54740
rect 86184 54684 86240 54740
rect 85812 54560 85868 54616
rect 85936 54560 85992 54616
rect 86060 54560 86116 54616
rect 86184 54560 86240 54616
rect 85812 54436 85868 54492
rect 85936 54436 85992 54492
rect 86060 54436 86116 54492
rect 86184 54436 86240 54492
rect 86612 53908 86668 53964
rect 86736 53908 86792 53964
rect 86860 53908 86916 53964
rect 86984 53908 87040 53964
rect 1930 53784 1986 53840
rect 2054 53784 2110 53840
rect 2178 53784 2234 53840
rect 2302 53784 2358 53840
rect 1930 53660 1986 53716
rect 2054 53660 2110 53716
rect 2178 53660 2234 53716
rect 2302 53660 2358 53716
rect 86612 53784 86668 53840
rect 86736 53784 86792 53840
rect 86860 53784 86916 53840
rect 86984 53784 87040 53840
rect 86612 53660 86668 53716
rect 86736 53660 86792 53716
rect 86860 53660 86916 53716
rect 86984 53660 87040 53716
rect 86612 53536 86668 53592
rect 86736 53536 86792 53592
rect 86860 53536 86916 53592
rect 86984 53536 87040 53592
rect 1130 53008 1186 53064
rect 1254 53008 1310 53064
rect 1378 53008 1434 53064
rect 1502 53008 1558 53064
rect 1130 52884 1186 52940
rect 1254 52884 1310 52940
rect 1378 52884 1434 52940
rect 1502 52884 1558 52940
rect 1130 52760 1186 52816
rect 1254 52760 1310 52816
rect 1378 52760 1434 52816
rect 1502 52760 1558 52816
rect 1130 52636 1186 52692
rect 1254 52636 1310 52692
rect 1378 52636 1434 52692
rect 1502 52636 1558 52692
rect 85812 53008 85868 53064
rect 85936 53008 85992 53064
rect 86060 53008 86116 53064
rect 86184 53008 86240 53064
rect 85812 52884 85868 52940
rect 85936 52884 85992 52940
rect 86060 52884 86116 52940
rect 86184 52884 86240 52940
rect 85812 52760 85868 52816
rect 85936 52760 85992 52816
rect 86060 52760 86116 52816
rect 86184 52760 86240 52816
rect 85812 52636 85868 52692
rect 85936 52636 85992 52692
rect 86060 52636 86116 52692
rect 86184 52636 86240 52692
rect 86612 52108 86668 52164
rect 86736 52108 86792 52164
rect 86860 52108 86916 52164
rect 86984 52108 87040 52164
rect 1930 51984 1986 52040
rect 2054 51984 2110 52040
rect 2178 51984 2234 52040
rect 2302 51984 2358 52040
rect 1930 51860 1986 51916
rect 2054 51860 2110 51916
rect 2178 51860 2234 51916
rect 2302 51860 2358 51916
rect 86612 51984 86668 52040
rect 86736 51984 86792 52040
rect 86860 51984 86916 52040
rect 86984 51984 87040 52040
rect 86612 51860 86668 51916
rect 86736 51860 86792 51916
rect 86860 51860 86916 51916
rect 86984 51860 87040 51916
rect 86612 51736 86668 51792
rect 86736 51736 86792 51792
rect 86860 51736 86916 51792
rect 86984 51736 87040 51792
rect 1130 51208 1186 51264
rect 1254 51208 1310 51264
rect 1378 51208 1434 51264
rect 1502 51208 1558 51264
rect 1130 51084 1186 51140
rect 1254 51084 1310 51140
rect 1378 51084 1434 51140
rect 1502 51084 1558 51140
rect 1130 50960 1186 51016
rect 1254 50960 1310 51016
rect 1378 50960 1434 51016
rect 1502 50960 1558 51016
rect 1130 50836 1186 50892
rect 1254 50836 1310 50892
rect 1378 50836 1434 50892
rect 1502 50836 1558 50892
rect 85812 51208 85868 51264
rect 85936 51208 85992 51264
rect 86060 51208 86116 51264
rect 86184 51208 86240 51264
rect 85812 51084 85868 51140
rect 85936 51084 85992 51140
rect 86060 51084 86116 51140
rect 86184 51084 86240 51140
rect 85812 50960 85868 51016
rect 85936 50960 85992 51016
rect 86060 50960 86116 51016
rect 86184 50960 86240 51016
rect 85812 50836 85868 50892
rect 85936 50836 85992 50892
rect 86060 50836 86116 50892
rect 86184 50836 86240 50892
rect 86612 50308 86668 50364
rect 86736 50308 86792 50364
rect 86860 50308 86916 50364
rect 86984 50308 87040 50364
rect 1930 50184 1986 50240
rect 2054 50184 2110 50240
rect 2178 50184 2234 50240
rect 2302 50184 2358 50240
rect 1930 50060 1986 50116
rect 2054 50060 2110 50116
rect 2178 50060 2234 50116
rect 2302 50060 2358 50116
rect 86612 50184 86668 50240
rect 86736 50184 86792 50240
rect 86860 50184 86916 50240
rect 86984 50184 87040 50240
rect 86612 50060 86668 50116
rect 86736 50060 86792 50116
rect 86860 50060 86916 50116
rect 86984 50060 87040 50116
rect 86612 49936 86668 49992
rect 86736 49936 86792 49992
rect 86860 49936 86916 49992
rect 86984 49936 87040 49992
rect 1130 49408 1186 49464
rect 1254 49408 1310 49464
rect 1378 49408 1434 49464
rect 1502 49408 1558 49464
rect 1130 49284 1186 49340
rect 1254 49284 1310 49340
rect 1378 49284 1434 49340
rect 1502 49284 1558 49340
rect 1130 49160 1186 49216
rect 1254 49160 1310 49216
rect 1378 49160 1434 49216
rect 1502 49160 1558 49216
rect 1130 49036 1186 49092
rect 1254 49036 1310 49092
rect 1378 49036 1434 49092
rect 1502 49036 1558 49092
rect 85812 49408 85868 49464
rect 85936 49408 85992 49464
rect 86060 49408 86116 49464
rect 86184 49408 86240 49464
rect 85812 49284 85868 49340
rect 85936 49284 85992 49340
rect 86060 49284 86116 49340
rect 86184 49284 86240 49340
rect 85812 49160 85868 49216
rect 85936 49160 85992 49216
rect 86060 49160 86116 49216
rect 86184 49160 86240 49216
rect 85812 49036 85868 49092
rect 85936 49036 85992 49092
rect 86060 49036 86116 49092
rect 86184 49036 86240 49092
rect 86612 48508 86668 48564
rect 86736 48508 86792 48564
rect 86860 48508 86916 48564
rect 86984 48508 87040 48564
rect 1930 48384 1986 48440
rect 2054 48384 2110 48440
rect 2178 48384 2234 48440
rect 2302 48384 2358 48440
rect 1930 48260 1986 48316
rect 2054 48260 2110 48316
rect 2178 48260 2234 48316
rect 2302 48260 2358 48316
rect 86612 48384 86668 48440
rect 86736 48384 86792 48440
rect 86860 48384 86916 48440
rect 86984 48384 87040 48440
rect 86612 48260 86668 48316
rect 86736 48260 86792 48316
rect 86860 48260 86916 48316
rect 86984 48260 87040 48316
rect 86612 48136 86668 48192
rect 86736 48136 86792 48192
rect 86860 48136 86916 48192
rect 86984 48136 87040 48192
rect 1130 47608 1186 47664
rect 1254 47608 1310 47664
rect 1378 47608 1434 47664
rect 1502 47608 1558 47664
rect 1130 47484 1186 47540
rect 1254 47484 1310 47540
rect 1378 47484 1434 47540
rect 1502 47484 1558 47540
rect 1130 47360 1186 47416
rect 1254 47360 1310 47416
rect 1378 47360 1434 47416
rect 1502 47360 1558 47416
rect 1130 47236 1186 47292
rect 1254 47236 1310 47292
rect 1378 47236 1434 47292
rect 1502 47236 1558 47292
rect 85812 47608 85868 47664
rect 85936 47608 85992 47664
rect 86060 47608 86116 47664
rect 86184 47608 86240 47664
rect 85812 47484 85868 47540
rect 85936 47484 85992 47540
rect 86060 47484 86116 47540
rect 86184 47484 86240 47540
rect 85812 47360 85868 47416
rect 85936 47360 85992 47416
rect 86060 47360 86116 47416
rect 86184 47360 86240 47416
rect 85812 47236 85868 47292
rect 85936 47236 85992 47292
rect 86060 47236 86116 47292
rect 86184 47236 86240 47292
rect 86612 46708 86668 46764
rect 86736 46708 86792 46764
rect 86860 46708 86916 46764
rect 86984 46708 87040 46764
rect 1930 46584 1986 46640
rect 2054 46584 2110 46640
rect 2178 46584 2234 46640
rect 2302 46584 2358 46640
rect 1930 46460 1986 46516
rect 2054 46460 2110 46516
rect 2178 46460 2234 46516
rect 2302 46460 2358 46516
rect 86612 46584 86668 46640
rect 86736 46584 86792 46640
rect 86860 46584 86916 46640
rect 86984 46584 87040 46640
rect 86612 46460 86668 46516
rect 86736 46460 86792 46516
rect 86860 46460 86916 46516
rect 86984 46460 87040 46516
rect 86612 46336 86668 46392
rect 86736 46336 86792 46392
rect 86860 46336 86916 46392
rect 86984 46336 87040 46392
rect 1130 45808 1186 45864
rect 1254 45808 1310 45864
rect 1378 45808 1434 45864
rect 1502 45808 1558 45864
rect 1130 45684 1186 45740
rect 1254 45684 1310 45740
rect 1378 45684 1434 45740
rect 1502 45684 1558 45740
rect 1130 45560 1186 45616
rect 1254 45560 1310 45616
rect 1378 45560 1434 45616
rect 1502 45560 1558 45616
rect 1130 45436 1186 45492
rect 1254 45436 1310 45492
rect 1378 45436 1434 45492
rect 1502 45436 1558 45492
rect 85812 45808 85868 45864
rect 85936 45808 85992 45864
rect 86060 45808 86116 45864
rect 86184 45808 86240 45864
rect 85812 45684 85868 45740
rect 85936 45684 85992 45740
rect 86060 45684 86116 45740
rect 86184 45684 86240 45740
rect 85812 45560 85868 45616
rect 85936 45560 85992 45616
rect 86060 45560 86116 45616
rect 86184 45560 86240 45616
rect 85812 45436 85868 45492
rect 85936 45436 85992 45492
rect 86060 45436 86116 45492
rect 86184 45436 86240 45492
rect 86612 44908 86668 44964
rect 86736 44908 86792 44964
rect 86860 44908 86916 44964
rect 86984 44908 87040 44964
rect 1930 44784 1986 44840
rect 2054 44784 2110 44840
rect 2178 44784 2234 44840
rect 2302 44784 2358 44840
rect 1930 44660 1986 44716
rect 2054 44660 2110 44716
rect 2178 44660 2234 44716
rect 2302 44660 2358 44716
rect 86612 44784 86668 44840
rect 86736 44784 86792 44840
rect 86860 44784 86916 44840
rect 86984 44784 87040 44840
rect 86612 44660 86668 44716
rect 86736 44660 86792 44716
rect 86860 44660 86916 44716
rect 86984 44660 87040 44716
rect 86612 44536 86668 44592
rect 86736 44536 86792 44592
rect 86860 44536 86916 44592
rect 86984 44536 87040 44592
rect 1130 44008 1186 44064
rect 1254 44008 1310 44064
rect 1378 44008 1434 44064
rect 1502 44008 1558 44064
rect 1130 43884 1186 43940
rect 1254 43884 1310 43940
rect 1378 43884 1434 43940
rect 1502 43884 1558 43940
rect 1130 43760 1186 43816
rect 1254 43760 1310 43816
rect 1378 43760 1434 43816
rect 1502 43760 1558 43816
rect 1130 43636 1186 43692
rect 1254 43636 1310 43692
rect 1378 43636 1434 43692
rect 1502 43636 1558 43692
rect 85812 44008 85868 44064
rect 85936 44008 85992 44064
rect 86060 44008 86116 44064
rect 86184 44008 86240 44064
rect 85812 43884 85868 43940
rect 85936 43884 85992 43940
rect 86060 43884 86116 43940
rect 86184 43884 86240 43940
rect 85812 43760 85868 43816
rect 85936 43760 85992 43816
rect 86060 43760 86116 43816
rect 86184 43760 86240 43816
rect 85812 43636 85868 43692
rect 85936 43636 85992 43692
rect 86060 43636 86116 43692
rect 86184 43636 86240 43692
rect 86612 43108 86668 43164
rect 86736 43108 86792 43164
rect 86860 43108 86916 43164
rect 86984 43108 87040 43164
rect 1930 42984 1986 43040
rect 2054 42984 2110 43040
rect 2178 42984 2234 43040
rect 2302 42984 2358 43040
rect 1930 42860 1986 42916
rect 2054 42860 2110 42916
rect 2178 42860 2234 42916
rect 2302 42860 2358 42916
rect 86612 42984 86668 43040
rect 86736 42984 86792 43040
rect 86860 42984 86916 43040
rect 86984 42984 87040 43040
rect 86612 42860 86668 42916
rect 86736 42860 86792 42916
rect 86860 42860 86916 42916
rect 86984 42860 87040 42916
rect 86612 42736 86668 42792
rect 86736 42736 86792 42792
rect 86860 42736 86916 42792
rect 86984 42736 87040 42792
rect 1130 42208 1186 42264
rect 1254 42208 1310 42264
rect 1378 42208 1434 42264
rect 1502 42208 1558 42264
rect 1130 42084 1186 42140
rect 1254 42084 1310 42140
rect 1378 42084 1434 42140
rect 1502 42084 1558 42140
rect 1130 41960 1186 42016
rect 1254 41960 1310 42016
rect 1378 41960 1434 42016
rect 1502 41960 1558 42016
rect 1130 41836 1186 41892
rect 1254 41836 1310 41892
rect 1378 41836 1434 41892
rect 1502 41836 1558 41892
rect 85812 42208 85868 42264
rect 85936 42208 85992 42264
rect 86060 42208 86116 42264
rect 86184 42208 86240 42264
rect 85812 42084 85868 42140
rect 85936 42084 85992 42140
rect 86060 42084 86116 42140
rect 86184 42084 86240 42140
rect 85812 41960 85868 42016
rect 85936 41960 85992 42016
rect 86060 41960 86116 42016
rect 86184 41960 86240 42016
rect 85812 41836 85868 41892
rect 85936 41836 85992 41892
rect 86060 41836 86116 41892
rect 86184 41836 86240 41892
rect 86612 41308 86668 41364
rect 86736 41308 86792 41364
rect 86860 41308 86916 41364
rect 86984 41308 87040 41364
rect 1930 41184 1986 41240
rect 2054 41184 2110 41240
rect 2178 41184 2234 41240
rect 2302 41184 2358 41240
rect 1930 41060 1986 41116
rect 2054 41060 2110 41116
rect 2178 41060 2234 41116
rect 2302 41060 2358 41116
rect 86612 41184 86668 41240
rect 86736 41184 86792 41240
rect 86860 41184 86916 41240
rect 86984 41184 87040 41240
rect 86612 41060 86668 41116
rect 86736 41060 86792 41116
rect 86860 41060 86916 41116
rect 86984 41060 87040 41116
rect 86612 40936 86668 40992
rect 86736 40936 86792 40992
rect 86860 40936 86916 40992
rect 86984 40936 87040 40992
rect 1130 40408 1186 40464
rect 1254 40408 1310 40464
rect 1378 40408 1434 40464
rect 1502 40408 1558 40464
rect 1130 40284 1186 40340
rect 1254 40284 1310 40340
rect 1378 40284 1434 40340
rect 1502 40284 1558 40340
rect 1130 40160 1186 40216
rect 1254 40160 1310 40216
rect 1378 40160 1434 40216
rect 1502 40160 1558 40216
rect 1130 40036 1186 40092
rect 1254 40036 1310 40092
rect 1378 40036 1434 40092
rect 1502 40036 1558 40092
rect 85812 40408 85868 40464
rect 85936 40408 85992 40464
rect 86060 40408 86116 40464
rect 86184 40408 86240 40464
rect 85812 40284 85868 40340
rect 85936 40284 85992 40340
rect 86060 40284 86116 40340
rect 86184 40284 86240 40340
rect 85812 40160 85868 40216
rect 85936 40160 85992 40216
rect 86060 40160 86116 40216
rect 86184 40160 86240 40216
rect 85812 40036 85868 40092
rect 85936 40036 85992 40092
rect 86060 40036 86116 40092
rect 86184 40036 86240 40092
rect 86612 39508 86668 39564
rect 86736 39508 86792 39564
rect 86860 39508 86916 39564
rect 86984 39508 87040 39564
rect 1930 39384 1986 39440
rect 2054 39384 2110 39440
rect 2178 39384 2234 39440
rect 2302 39384 2358 39440
rect 1930 39260 1986 39316
rect 2054 39260 2110 39316
rect 2178 39260 2234 39316
rect 2302 39260 2358 39316
rect 86612 39384 86668 39440
rect 86736 39384 86792 39440
rect 86860 39384 86916 39440
rect 86984 39384 87040 39440
rect 86612 39260 86668 39316
rect 86736 39260 86792 39316
rect 86860 39260 86916 39316
rect 86984 39260 87040 39316
rect 86612 39136 86668 39192
rect 86736 39136 86792 39192
rect 86860 39136 86916 39192
rect 86984 39136 87040 39192
rect 1130 38608 1186 38664
rect 1254 38608 1310 38664
rect 1378 38608 1434 38664
rect 1502 38608 1558 38664
rect 1130 38484 1186 38540
rect 1254 38484 1310 38540
rect 1378 38484 1434 38540
rect 1502 38484 1558 38540
rect 1130 38360 1186 38416
rect 1254 38360 1310 38416
rect 1378 38360 1434 38416
rect 1502 38360 1558 38416
rect 1130 38236 1186 38292
rect 1254 38236 1310 38292
rect 1378 38236 1434 38292
rect 1502 38236 1558 38292
rect 85812 38608 85868 38664
rect 85936 38608 85992 38664
rect 86060 38608 86116 38664
rect 86184 38608 86240 38664
rect 85812 38484 85868 38540
rect 85936 38484 85992 38540
rect 86060 38484 86116 38540
rect 86184 38484 86240 38540
rect 85812 38360 85868 38416
rect 85936 38360 85992 38416
rect 86060 38360 86116 38416
rect 86184 38360 86240 38416
rect 85812 38236 85868 38292
rect 85936 38236 85992 38292
rect 86060 38236 86116 38292
rect 86184 38236 86240 38292
rect 86612 37708 86668 37764
rect 86736 37708 86792 37764
rect 86860 37708 86916 37764
rect 86984 37708 87040 37764
rect 1930 37584 1986 37640
rect 2054 37584 2110 37640
rect 2178 37584 2234 37640
rect 2302 37584 2358 37640
rect 1930 37460 1986 37516
rect 2054 37460 2110 37516
rect 2178 37460 2234 37516
rect 2302 37460 2358 37516
rect 86612 37584 86668 37640
rect 86736 37584 86792 37640
rect 86860 37584 86916 37640
rect 86984 37584 87040 37640
rect 86612 37460 86668 37516
rect 86736 37460 86792 37516
rect 86860 37460 86916 37516
rect 86984 37460 87040 37516
rect 86612 37336 86668 37392
rect 86736 37336 86792 37392
rect 86860 37336 86916 37392
rect 86984 37336 87040 37392
rect 1130 36808 1186 36864
rect 1254 36808 1310 36864
rect 1378 36808 1434 36864
rect 1502 36808 1558 36864
rect 1130 36684 1186 36740
rect 1254 36684 1310 36740
rect 1378 36684 1434 36740
rect 1502 36684 1558 36740
rect 1130 36560 1186 36616
rect 1254 36560 1310 36616
rect 1378 36560 1434 36616
rect 1502 36560 1558 36616
rect 1130 36436 1186 36492
rect 1254 36436 1310 36492
rect 1378 36436 1434 36492
rect 1502 36436 1558 36492
rect 85812 36808 85868 36864
rect 85936 36808 85992 36864
rect 86060 36808 86116 36864
rect 86184 36808 86240 36864
rect 85812 36684 85868 36740
rect 85936 36684 85992 36740
rect 86060 36684 86116 36740
rect 86184 36684 86240 36740
rect 85812 36560 85868 36616
rect 85936 36560 85992 36616
rect 86060 36560 86116 36616
rect 86184 36560 86240 36616
rect 85812 36436 85868 36492
rect 85936 36436 85992 36492
rect 86060 36436 86116 36492
rect 86184 36436 86240 36492
rect 86612 35908 86668 35964
rect 86736 35908 86792 35964
rect 86860 35908 86916 35964
rect 86984 35908 87040 35964
rect 1930 35784 1986 35840
rect 2054 35784 2110 35840
rect 2178 35784 2234 35840
rect 2302 35784 2358 35840
rect 1930 35660 1986 35716
rect 2054 35660 2110 35716
rect 2178 35660 2234 35716
rect 2302 35660 2358 35716
rect 86612 35784 86668 35840
rect 86736 35784 86792 35840
rect 86860 35784 86916 35840
rect 86984 35784 87040 35840
rect 86612 35660 86668 35716
rect 86736 35660 86792 35716
rect 86860 35660 86916 35716
rect 86984 35660 87040 35716
rect 86612 35536 86668 35592
rect 86736 35536 86792 35592
rect 86860 35536 86916 35592
rect 86984 35536 87040 35592
rect 1130 35008 1186 35064
rect 1254 35008 1310 35064
rect 1378 35008 1434 35064
rect 1502 35008 1558 35064
rect 1130 34884 1186 34940
rect 1254 34884 1310 34940
rect 1378 34884 1434 34940
rect 1502 34884 1558 34940
rect 1130 34760 1186 34816
rect 1254 34760 1310 34816
rect 1378 34760 1434 34816
rect 1502 34760 1558 34816
rect 1130 34636 1186 34692
rect 1254 34636 1310 34692
rect 1378 34636 1434 34692
rect 1502 34636 1558 34692
rect 85812 35008 85868 35064
rect 85936 35008 85992 35064
rect 86060 35008 86116 35064
rect 86184 35008 86240 35064
rect 85812 34884 85868 34940
rect 85936 34884 85992 34940
rect 86060 34884 86116 34940
rect 86184 34884 86240 34940
rect 85812 34760 85868 34816
rect 85936 34760 85992 34816
rect 86060 34760 86116 34816
rect 86184 34760 86240 34816
rect 85812 34636 85868 34692
rect 85936 34636 85992 34692
rect 86060 34636 86116 34692
rect 86184 34636 86240 34692
rect 86612 34108 86668 34164
rect 86736 34108 86792 34164
rect 86860 34108 86916 34164
rect 86984 34108 87040 34164
rect 1930 33984 1986 34040
rect 2054 33984 2110 34040
rect 2178 33984 2234 34040
rect 2302 33984 2358 34040
rect 1930 33860 1986 33916
rect 2054 33860 2110 33916
rect 2178 33860 2234 33916
rect 2302 33860 2358 33916
rect 86612 33984 86668 34040
rect 86736 33984 86792 34040
rect 86860 33984 86916 34040
rect 86984 33984 87040 34040
rect 86612 33860 86668 33916
rect 86736 33860 86792 33916
rect 86860 33860 86916 33916
rect 86984 33860 87040 33916
rect 86612 33736 86668 33792
rect 86736 33736 86792 33792
rect 86860 33736 86916 33792
rect 86984 33736 87040 33792
rect 1130 33208 1186 33264
rect 1254 33208 1310 33264
rect 1378 33208 1434 33264
rect 1502 33208 1558 33264
rect 1130 33084 1186 33140
rect 1254 33084 1310 33140
rect 1378 33084 1434 33140
rect 1502 33084 1558 33140
rect 1130 32960 1186 33016
rect 1254 32960 1310 33016
rect 1378 32960 1434 33016
rect 1502 32960 1558 33016
rect 1130 32836 1186 32892
rect 1254 32836 1310 32892
rect 1378 32836 1434 32892
rect 1502 32836 1558 32892
rect 85812 33208 85868 33264
rect 85936 33208 85992 33264
rect 86060 33208 86116 33264
rect 86184 33208 86240 33264
rect 85812 33084 85868 33140
rect 85936 33084 85992 33140
rect 86060 33084 86116 33140
rect 86184 33084 86240 33140
rect 85812 32960 85868 33016
rect 85936 32960 85992 33016
rect 86060 32960 86116 33016
rect 86184 32960 86240 33016
rect 85812 32836 85868 32892
rect 85936 32836 85992 32892
rect 86060 32836 86116 32892
rect 86184 32836 86240 32892
rect 86612 32308 86668 32364
rect 86736 32308 86792 32364
rect 86860 32308 86916 32364
rect 86984 32308 87040 32364
rect 1930 32184 1986 32240
rect 2054 32184 2110 32240
rect 2178 32184 2234 32240
rect 2302 32184 2358 32240
rect 1930 32060 1986 32116
rect 2054 32060 2110 32116
rect 2178 32060 2234 32116
rect 2302 32060 2358 32116
rect 86612 32184 86668 32240
rect 86736 32184 86792 32240
rect 86860 32184 86916 32240
rect 86984 32184 87040 32240
rect 86612 32060 86668 32116
rect 86736 32060 86792 32116
rect 86860 32060 86916 32116
rect 86984 32060 87040 32116
rect 86612 31936 86668 31992
rect 86736 31936 86792 31992
rect 86860 31936 86916 31992
rect 86984 31936 87040 31992
rect 1130 31408 1186 31464
rect 1254 31408 1310 31464
rect 1378 31408 1434 31464
rect 1502 31408 1558 31464
rect 1130 31284 1186 31340
rect 1254 31284 1310 31340
rect 1378 31284 1434 31340
rect 1502 31284 1558 31340
rect 1130 31160 1186 31216
rect 1254 31160 1310 31216
rect 1378 31160 1434 31216
rect 1502 31160 1558 31216
rect 1130 31036 1186 31092
rect 1254 31036 1310 31092
rect 1378 31036 1434 31092
rect 1502 31036 1558 31092
rect 85812 31408 85868 31464
rect 85936 31408 85992 31464
rect 86060 31408 86116 31464
rect 86184 31408 86240 31464
rect 85812 31284 85868 31340
rect 85936 31284 85992 31340
rect 86060 31284 86116 31340
rect 86184 31284 86240 31340
rect 85812 31160 85868 31216
rect 85936 31160 85992 31216
rect 86060 31160 86116 31216
rect 86184 31160 86240 31216
rect 85812 31036 85868 31092
rect 85936 31036 85992 31092
rect 86060 31036 86116 31092
rect 86184 31036 86240 31092
rect 86612 30508 86668 30564
rect 86736 30508 86792 30564
rect 86860 30508 86916 30564
rect 86984 30508 87040 30564
rect 1930 30384 1986 30440
rect 2054 30384 2110 30440
rect 2178 30384 2234 30440
rect 2302 30384 2358 30440
rect 1930 30260 1986 30316
rect 2054 30260 2110 30316
rect 2178 30260 2234 30316
rect 2302 30260 2358 30316
rect 86612 30384 86668 30440
rect 86736 30384 86792 30440
rect 86860 30384 86916 30440
rect 86984 30384 87040 30440
rect 86612 30260 86668 30316
rect 86736 30260 86792 30316
rect 86860 30260 86916 30316
rect 86984 30260 87040 30316
rect 86612 30136 86668 30192
rect 86736 30136 86792 30192
rect 86860 30136 86916 30192
rect 86984 30136 87040 30192
rect 1130 29608 1186 29664
rect 1254 29608 1310 29664
rect 1378 29608 1434 29664
rect 1502 29608 1558 29664
rect 1130 29484 1186 29540
rect 1254 29484 1310 29540
rect 1378 29484 1434 29540
rect 1502 29484 1558 29540
rect 1130 29360 1186 29416
rect 1254 29360 1310 29416
rect 1378 29360 1434 29416
rect 1502 29360 1558 29416
rect 1130 29236 1186 29292
rect 1254 29236 1310 29292
rect 1378 29236 1434 29292
rect 1502 29236 1558 29292
rect 85812 29608 85868 29664
rect 85936 29608 85992 29664
rect 86060 29608 86116 29664
rect 86184 29608 86240 29664
rect 85812 29484 85868 29540
rect 85936 29484 85992 29540
rect 86060 29484 86116 29540
rect 86184 29484 86240 29540
rect 85812 29360 85868 29416
rect 85936 29360 85992 29416
rect 86060 29360 86116 29416
rect 86184 29360 86240 29416
rect 85812 29236 85868 29292
rect 85936 29236 85992 29292
rect 86060 29236 86116 29292
rect 86184 29236 86240 29292
rect 86612 28708 86668 28764
rect 86736 28708 86792 28764
rect 86860 28708 86916 28764
rect 86984 28708 87040 28764
rect 1930 28584 1986 28640
rect 2054 28584 2110 28640
rect 2178 28584 2234 28640
rect 2302 28584 2358 28640
rect 1930 28460 1986 28516
rect 2054 28460 2110 28516
rect 2178 28460 2234 28516
rect 2302 28460 2358 28516
rect 86612 28584 86668 28640
rect 86736 28584 86792 28640
rect 86860 28584 86916 28640
rect 86984 28584 87040 28640
rect 86612 28460 86668 28516
rect 86736 28460 86792 28516
rect 86860 28460 86916 28516
rect 86984 28460 87040 28516
rect 86612 28336 86668 28392
rect 86736 28336 86792 28392
rect 86860 28336 86916 28392
rect 86984 28336 87040 28392
rect 1130 27808 1186 27864
rect 1254 27808 1310 27864
rect 1378 27808 1434 27864
rect 1502 27808 1558 27864
rect 1130 27684 1186 27740
rect 1254 27684 1310 27740
rect 1378 27684 1434 27740
rect 1502 27684 1558 27740
rect 1130 27560 1186 27616
rect 1254 27560 1310 27616
rect 1378 27560 1434 27616
rect 1502 27560 1558 27616
rect 1130 27436 1186 27492
rect 1254 27436 1310 27492
rect 1378 27436 1434 27492
rect 1502 27436 1558 27492
rect 85812 27808 85868 27864
rect 85936 27808 85992 27864
rect 86060 27808 86116 27864
rect 86184 27808 86240 27864
rect 85812 27684 85868 27740
rect 85936 27684 85992 27740
rect 86060 27684 86116 27740
rect 86184 27684 86240 27740
rect 85812 27560 85868 27616
rect 85936 27560 85992 27616
rect 86060 27560 86116 27616
rect 86184 27560 86240 27616
rect 85812 27436 85868 27492
rect 85936 27436 85992 27492
rect 86060 27436 86116 27492
rect 86184 27436 86240 27492
rect 86612 26908 86668 26964
rect 86736 26908 86792 26964
rect 86860 26908 86916 26964
rect 86984 26908 87040 26964
rect 1930 26784 1986 26840
rect 2054 26784 2110 26840
rect 2178 26784 2234 26840
rect 2302 26784 2358 26840
rect 1930 26660 1986 26716
rect 2054 26660 2110 26716
rect 2178 26660 2234 26716
rect 2302 26660 2358 26716
rect 86612 26784 86668 26840
rect 86736 26784 86792 26840
rect 86860 26784 86916 26840
rect 86984 26784 87040 26840
rect 86612 26660 86668 26716
rect 86736 26660 86792 26716
rect 86860 26660 86916 26716
rect 86984 26660 87040 26716
rect 86612 26536 86668 26592
rect 86736 26536 86792 26592
rect 86860 26536 86916 26592
rect 86984 26536 87040 26592
rect 1130 26008 1186 26064
rect 1254 26008 1310 26064
rect 1378 26008 1434 26064
rect 1502 26008 1558 26064
rect 1130 25884 1186 25940
rect 1254 25884 1310 25940
rect 1378 25884 1434 25940
rect 1502 25884 1558 25940
rect 1130 25760 1186 25816
rect 1254 25760 1310 25816
rect 1378 25760 1434 25816
rect 1502 25760 1558 25816
rect 1130 25636 1186 25692
rect 1254 25636 1310 25692
rect 1378 25636 1434 25692
rect 1502 25636 1558 25692
rect 85812 26008 85868 26064
rect 85936 26008 85992 26064
rect 86060 26008 86116 26064
rect 86184 26008 86240 26064
rect 85812 25884 85868 25940
rect 85936 25884 85992 25940
rect 86060 25884 86116 25940
rect 86184 25884 86240 25940
rect 85812 25760 85868 25816
rect 85936 25760 85992 25816
rect 86060 25760 86116 25816
rect 86184 25760 86240 25816
rect 85812 25636 85868 25692
rect 85936 25636 85992 25692
rect 86060 25636 86116 25692
rect 86184 25636 86240 25692
rect 86612 25108 86668 25164
rect 86736 25108 86792 25164
rect 86860 25108 86916 25164
rect 86984 25108 87040 25164
rect 1930 24984 1986 25040
rect 2054 24984 2110 25040
rect 2178 24984 2234 25040
rect 2302 24984 2358 25040
rect 1930 24860 1986 24916
rect 2054 24860 2110 24916
rect 2178 24860 2234 24916
rect 2302 24860 2358 24916
rect 86612 24984 86668 25040
rect 86736 24984 86792 25040
rect 86860 24984 86916 25040
rect 86984 24984 87040 25040
rect 86612 24860 86668 24916
rect 86736 24860 86792 24916
rect 86860 24860 86916 24916
rect 86984 24860 87040 24916
rect 86612 24736 86668 24792
rect 86736 24736 86792 24792
rect 86860 24736 86916 24792
rect 86984 24736 87040 24792
rect 1130 24208 1186 24264
rect 1254 24208 1310 24264
rect 1378 24208 1434 24264
rect 1502 24208 1558 24264
rect 1130 24084 1186 24140
rect 1254 24084 1310 24140
rect 1378 24084 1434 24140
rect 1502 24084 1558 24140
rect 1130 23960 1186 24016
rect 1254 23960 1310 24016
rect 1378 23960 1434 24016
rect 1502 23960 1558 24016
rect 1130 23836 1186 23892
rect 1254 23836 1310 23892
rect 1378 23836 1434 23892
rect 1502 23836 1558 23892
rect 85812 24208 85868 24264
rect 85936 24208 85992 24264
rect 86060 24208 86116 24264
rect 86184 24208 86240 24264
rect 85812 24084 85868 24140
rect 85936 24084 85992 24140
rect 86060 24084 86116 24140
rect 86184 24084 86240 24140
rect 85812 23960 85868 24016
rect 85936 23960 85992 24016
rect 86060 23960 86116 24016
rect 86184 23960 86240 24016
rect 85812 23836 85868 23892
rect 85936 23836 85992 23892
rect 86060 23836 86116 23892
rect 86184 23836 86240 23892
rect 86612 23308 86668 23364
rect 86736 23308 86792 23364
rect 86860 23308 86916 23364
rect 86984 23308 87040 23364
rect 1930 23184 1986 23240
rect 2054 23184 2110 23240
rect 2178 23184 2234 23240
rect 2302 23184 2358 23240
rect 1930 23060 1986 23116
rect 2054 23060 2110 23116
rect 2178 23060 2234 23116
rect 2302 23060 2358 23116
rect 86612 23184 86668 23240
rect 86736 23184 86792 23240
rect 86860 23184 86916 23240
rect 86984 23184 87040 23240
rect 86612 23060 86668 23116
rect 86736 23060 86792 23116
rect 86860 23060 86916 23116
rect 86984 23060 87040 23116
rect 86612 22936 86668 22992
rect 86736 22936 86792 22992
rect 86860 22936 86916 22992
rect 86984 22936 87040 22992
rect 1130 22408 1186 22464
rect 1254 22408 1310 22464
rect 1378 22408 1434 22464
rect 1502 22408 1558 22464
rect 1130 22284 1186 22340
rect 1254 22284 1310 22340
rect 1378 22284 1434 22340
rect 1502 22284 1558 22340
rect 1130 22160 1186 22216
rect 1254 22160 1310 22216
rect 1378 22160 1434 22216
rect 1502 22160 1558 22216
rect 1130 22036 1186 22092
rect 1254 22036 1310 22092
rect 1378 22036 1434 22092
rect 1502 22036 1558 22092
rect 85812 22408 85868 22464
rect 85936 22408 85992 22464
rect 86060 22408 86116 22464
rect 86184 22408 86240 22464
rect 85812 22284 85868 22340
rect 85936 22284 85992 22340
rect 86060 22284 86116 22340
rect 86184 22284 86240 22340
rect 85812 22160 85868 22216
rect 85936 22160 85992 22216
rect 86060 22160 86116 22216
rect 86184 22160 86240 22216
rect 85812 22036 85868 22092
rect 85936 22036 85992 22092
rect 86060 22036 86116 22092
rect 86184 22036 86240 22092
rect 86612 21508 86668 21564
rect 86736 21508 86792 21564
rect 86860 21508 86916 21564
rect 86984 21508 87040 21564
rect 1930 21384 1986 21440
rect 2054 21384 2110 21440
rect 2178 21384 2234 21440
rect 2302 21384 2358 21440
rect 1930 21260 1986 21316
rect 2054 21260 2110 21316
rect 2178 21260 2234 21316
rect 2302 21260 2358 21316
rect 86612 21384 86668 21440
rect 86736 21384 86792 21440
rect 86860 21384 86916 21440
rect 86984 21384 87040 21440
rect 86612 21260 86668 21316
rect 86736 21260 86792 21316
rect 86860 21260 86916 21316
rect 86984 21260 87040 21316
rect 86612 21136 86668 21192
rect 86736 21136 86792 21192
rect 86860 21136 86916 21192
rect 86984 21136 87040 21192
rect 1130 20608 1186 20664
rect 1254 20608 1310 20664
rect 1378 20608 1434 20664
rect 1502 20608 1558 20664
rect 1130 20484 1186 20540
rect 1254 20484 1310 20540
rect 1378 20484 1434 20540
rect 1502 20484 1558 20540
rect 1130 20360 1186 20416
rect 1254 20360 1310 20416
rect 1378 20360 1434 20416
rect 1502 20360 1558 20416
rect 1130 20236 1186 20292
rect 1254 20236 1310 20292
rect 1378 20236 1434 20292
rect 1502 20236 1558 20292
rect 85812 20608 85868 20664
rect 85936 20608 85992 20664
rect 86060 20608 86116 20664
rect 86184 20608 86240 20664
rect 85812 20484 85868 20540
rect 85936 20484 85992 20540
rect 86060 20484 86116 20540
rect 86184 20484 86240 20540
rect 85812 20360 85868 20416
rect 85936 20360 85992 20416
rect 86060 20360 86116 20416
rect 86184 20360 86240 20416
rect 85812 20236 85868 20292
rect 85936 20236 85992 20292
rect 86060 20236 86116 20292
rect 86184 20236 86240 20292
rect 86612 19708 86668 19764
rect 86736 19708 86792 19764
rect 86860 19708 86916 19764
rect 86984 19708 87040 19764
rect 1930 19584 1986 19640
rect 2054 19584 2110 19640
rect 2178 19584 2234 19640
rect 2302 19584 2358 19640
rect 1930 19460 1986 19516
rect 2054 19460 2110 19516
rect 2178 19460 2234 19516
rect 2302 19460 2358 19516
rect 86612 19584 86668 19640
rect 86736 19584 86792 19640
rect 86860 19584 86916 19640
rect 86984 19584 87040 19640
rect 86612 19460 86668 19516
rect 86736 19460 86792 19516
rect 86860 19460 86916 19516
rect 86984 19460 87040 19516
rect 86612 19336 86668 19392
rect 86736 19336 86792 19392
rect 86860 19336 86916 19392
rect 86984 19336 87040 19392
rect 1130 18808 1186 18864
rect 1254 18808 1310 18864
rect 1378 18808 1434 18864
rect 1502 18808 1558 18864
rect 1130 18684 1186 18740
rect 1254 18684 1310 18740
rect 1378 18684 1434 18740
rect 1502 18684 1558 18740
rect 1130 18560 1186 18616
rect 1254 18560 1310 18616
rect 1378 18560 1434 18616
rect 1502 18560 1558 18616
rect 1130 18436 1186 18492
rect 1254 18436 1310 18492
rect 1378 18436 1434 18492
rect 1502 18436 1558 18492
rect 85812 18808 85868 18864
rect 85936 18808 85992 18864
rect 86060 18808 86116 18864
rect 86184 18808 86240 18864
rect 85812 18684 85868 18740
rect 85936 18684 85992 18740
rect 86060 18684 86116 18740
rect 86184 18684 86240 18740
rect 85812 18560 85868 18616
rect 85936 18560 85992 18616
rect 86060 18560 86116 18616
rect 86184 18560 86240 18616
rect 85812 18436 85868 18492
rect 85936 18436 85992 18492
rect 86060 18436 86116 18492
rect 86184 18436 86240 18492
rect 86612 17908 86668 17964
rect 86736 17908 86792 17964
rect 86860 17908 86916 17964
rect 86984 17908 87040 17964
rect 1930 17784 1986 17840
rect 2054 17784 2110 17840
rect 2178 17784 2234 17840
rect 2302 17784 2358 17840
rect 1930 17660 1986 17716
rect 2054 17660 2110 17716
rect 2178 17660 2234 17716
rect 2302 17660 2358 17716
rect 86612 17784 86668 17840
rect 86736 17784 86792 17840
rect 86860 17784 86916 17840
rect 86984 17784 87040 17840
rect 86612 17660 86668 17716
rect 86736 17660 86792 17716
rect 86860 17660 86916 17716
rect 86984 17660 87040 17716
rect 86612 17536 86668 17592
rect 86736 17536 86792 17592
rect 86860 17536 86916 17592
rect 86984 17536 87040 17592
rect 1130 17008 1186 17064
rect 1254 17008 1310 17064
rect 1378 17008 1434 17064
rect 1502 17008 1558 17064
rect 1130 16884 1186 16940
rect 1254 16884 1310 16940
rect 1378 16884 1434 16940
rect 1502 16884 1558 16940
rect 1130 16760 1186 16816
rect 1254 16760 1310 16816
rect 1378 16760 1434 16816
rect 1502 16760 1558 16816
rect 1130 16636 1186 16692
rect 1254 16636 1310 16692
rect 1378 16636 1434 16692
rect 1502 16636 1558 16692
rect 85812 17008 85868 17064
rect 85936 17008 85992 17064
rect 86060 17008 86116 17064
rect 86184 17008 86240 17064
rect 85812 16884 85868 16940
rect 85936 16884 85992 16940
rect 86060 16884 86116 16940
rect 86184 16884 86240 16940
rect 85812 16760 85868 16816
rect 85936 16760 85992 16816
rect 86060 16760 86116 16816
rect 86184 16760 86240 16816
rect 85812 16636 85868 16692
rect 85936 16636 85992 16692
rect 86060 16636 86116 16692
rect 86184 16636 86240 16692
rect 86612 16108 86668 16164
rect 86736 16108 86792 16164
rect 86860 16108 86916 16164
rect 86984 16108 87040 16164
rect 1930 15984 1986 16040
rect 2054 15984 2110 16040
rect 2178 15984 2234 16040
rect 2302 15984 2358 16040
rect 1930 15860 1986 15916
rect 2054 15860 2110 15916
rect 2178 15860 2234 15916
rect 2302 15860 2358 15916
rect 86612 15984 86668 16040
rect 86736 15984 86792 16040
rect 86860 15984 86916 16040
rect 86984 15984 87040 16040
rect 86612 15860 86668 15916
rect 86736 15860 86792 15916
rect 86860 15860 86916 15916
rect 86984 15860 87040 15916
rect 86612 15736 86668 15792
rect 86736 15736 86792 15792
rect 86860 15736 86916 15792
rect 86984 15736 87040 15792
rect 1130 15208 1186 15264
rect 1254 15208 1310 15264
rect 1378 15208 1434 15264
rect 1502 15208 1558 15264
rect 1130 15084 1186 15140
rect 1254 15084 1310 15140
rect 1378 15084 1434 15140
rect 1502 15084 1558 15140
rect 1130 14960 1186 15016
rect 1254 14960 1310 15016
rect 1378 14960 1434 15016
rect 1502 14960 1558 15016
rect 1130 14836 1186 14892
rect 1254 14836 1310 14892
rect 1378 14836 1434 14892
rect 1502 14836 1558 14892
rect 85812 15208 85868 15264
rect 85936 15208 85992 15264
rect 86060 15208 86116 15264
rect 86184 15208 86240 15264
rect 85812 15084 85868 15140
rect 85936 15084 85992 15140
rect 86060 15084 86116 15140
rect 86184 15084 86240 15140
rect 85812 14960 85868 15016
rect 85936 14960 85992 15016
rect 86060 14960 86116 15016
rect 86184 14960 86240 15016
rect 85812 14836 85868 14892
rect 85936 14836 85992 14892
rect 86060 14836 86116 14892
rect 86184 14836 86240 14892
rect 86612 14308 86668 14364
rect 86736 14308 86792 14364
rect 86860 14308 86916 14364
rect 86984 14308 87040 14364
rect 1930 14184 1986 14240
rect 2054 14184 2110 14240
rect 2178 14184 2234 14240
rect 2302 14184 2358 14240
rect 1930 14060 1986 14116
rect 2054 14060 2110 14116
rect 2178 14060 2234 14116
rect 2302 14060 2358 14116
rect 86612 14184 86668 14240
rect 86736 14184 86792 14240
rect 86860 14184 86916 14240
rect 86984 14184 87040 14240
rect 86612 14060 86668 14116
rect 86736 14060 86792 14116
rect 86860 14060 86916 14116
rect 86984 14060 87040 14116
rect 86612 13936 86668 13992
rect 86736 13936 86792 13992
rect 86860 13936 86916 13992
rect 86984 13936 87040 13992
rect 1130 13408 1186 13464
rect 1254 13408 1310 13464
rect 1378 13408 1434 13464
rect 1502 13408 1558 13464
rect 1130 13284 1186 13340
rect 1254 13284 1310 13340
rect 1378 13284 1434 13340
rect 1502 13284 1558 13340
rect 1130 13160 1186 13216
rect 1254 13160 1310 13216
rect 1378 13160 1434 13216
rect 1502 13160 1558 13216
rect 1130 13036 1186 13092
rect 1254 13036 1310 13092
rect 1378 13036 1434 13092
rect 1502 13036 1558 13092
rect 85812 13408 85868 13464
rect 85936 13408 85992 13464
rect 86060 13408 86116 13464
rect 86184 13408 86240 13464
rect 85812 13284 85868 13340
rect 85936 13284 85992 13340
rect 86060 13284 86116 13340
rect 86184 13284 86240 13340
rect 85812 13160 85868 13216
rect 85936 13160 85992 13216
rect 86060 13160 86116 13216
rect 86184 13160 86240 13216
rect 85812 13036 85868 13092
rect 85936 13036 85992 13092
rect 86060 13036 86116 13092
rect 86184 13036 86240 13092
rect 86612 12508 86668 12564
rect 86736 12508 86792 12564
rect 86860 12508 86916 12564
rect 86984 12508 87040 12564
rect 1930 12384 1986 12440
rect 2054 12384 2110 12440
rect 2178 12384 2234 12440
rect 2302 12384 2358 12440
rect 1930 12260 1986 12316
rect 2054 12260 2110 12316
rect 2178 12260 2234 12316
rect 2302 12260 2358 12316
rect 86612 12384 86668 12440
rect 86736 12384 86792 12440
rect 86860 12384 86916 12440
rect 86984 12384 87040 12440
rect 86612 12260 86668 12316
rect 86736 12260 86792 12316
rect 86860 12260 86916 12316
rect 86984 12260 87040 12316
rect 86612 12136 86668 12192
rect 86736 12136 86792 12192
rect 86860 12136 86916 12192
rect 86984 12136 87040 12192
rect 1130 11608 1186 11664
rect 1254 11608 1310 11664
rect 1378 11608 1434 11664
rect 1502 11608 1558 11664
rect 1130 11484 1186 11540
rect 1254 11484 1310 11540
rect 1378 11484 1434 11540
rect 1502 11484 1558 11540
rect 1130 11360 1186 11416
rect 1254 11360 1310 11416
rect 1378 11360 1434 11416
rect 1502 11360 1558 11416
rect 1130 11236 1186 11292
rect 1254 11236 1310 11292
rect 1378 11236 1434 11292
rect 1502 11236 1558 11292
rect 85812 11608 85868 11664
rect 85936 11608 85992 11664
rect 86060 11608 86116 11664
rect 86184 11608 86240 11664
rect 85812 11484 85868 11540
rect 85936 11484 85992 11540
rect 86060 11484 86116 11540
rect 86184 11484 86240 11540
rect 85812 11360 85868 11416
rect 85936 11360 85992 11416
rect 86060 11360 86116 11416
rect 86184 11360 86240 11416
rect 85812 11236 85868 11292
rect 85936 11236 85992 11292
rect 86060 11236 86116 11292
rect 86184 11236 86240 11292
rect 86612 10708 86668 10764
rect 86736 10708 86792 10764
rect 86860 10708 86916 10764
rect 86984 10708 87040 10764
rect 1930 10584 1986 10640
rect 2054 10584 2110 10640
rect 2178 10584 2234 10640
rect 2302 10584 2358 10640
rect 1930 10460 1986 10516
rect 2054 10460 2110 10516
rect 2178 10460 2234 10516
rect 2302 10460 2358 10516
rect 86612 10584 86668 10640
rect 86736 10584 86792 10640
rect 86860 10584 86916 10640
rect 86984 10584 87040 10640
rect 86612 10460 86668 10516
rect 86736 10460 86792 10516
rect 86860 10460 86916 10516
rect 86984 10460 87040 10516
rect 86612 10336 86668 10392
rect 86736 10336 86792 10392
rect 86860 10336 86916 10392
rect 86984 10336 87040 10392
rect 1130 9808 1186 9864
rect 1254 9808 1310 9864
rect 1378 9808 1434 9864
rect 1502 9808 1558 9864
rect 1130 9684 1186 9740
rect 1254 9684 1310 9740
rect 1378 9684 1434 9740
rect 1502 9684 1558 9740
rect 1130 9560 1186 9616
rect 1254 9560 1310 9616
rect 1378 9560 1434 9616
rect 1502 9560 1558 9616
rect 1130 9436 1186 9492
rect 1254 9436 1310 9492
rect 1378 9436 1434 9492
rect 1502 9436 1558 9492
rect 85812 9808 85868 9864
rect 85936 9808 85992 9864
rect 86060 9808 86116 9864
rect 86184 9808 86240 9864
rect 85812 9684 85868 9740
rect 85936 9684 85992 9740
rect 86060 9684 86116 9740
rect 86184 9684 86240 9740
rect 85812 9560 85868 9616
rect 85936 9560 85992 9616
rect 86060 9560 86116 9616
rect 86184 9560 86240 9616
rect 85812 9436 85868 9492
rect 85936 9436 85992 9492
rect 86060 9436 86116 9492
rect 86184 9436 86240 9492
rect 86612 8908 86668 8964
rect 86736 8908 86792 8964
rect 86860 8908 86916 8964
rect 86984 8908 87040 8964
rect 1930 8784 1986 8840
rect 2054 8784 2110 8840
rect 2178 8784 2234 8840
rect 2302 8784 2358 8840
rect 1930 8660 1986 8716
rect 2054 8660 2110 8716
rect 2178 8660 2234 8716
rect 2302 8660 2358 8716
rect 86612 8784 86668 8840
rect 86736 8784 86792 8840
rect 86860 8784 86916 8840
rect 86984 8784 87040 8840
rect 86612 8660 86668 8716
rect 86736 8660 86792 8716
rect 86860 8660 86916 8716
rect 86984 8660 87040 8716
rect 86612 8536 86668 8592
rect 86736 8536 86792 8592
rect 86860 8536 86916 8592
rect 86984 8536 87040 8592
rect 1130 8008 1186 8064
rect 1254 8008 1310 8064
rect 1378 8008 1434 8064
rect 1502 8008 1558 8064
rect 1130 7884 1186 7940
rect 1254 7884 1310 7940
rect 1378 7884 1434 7940
rect 1502 7884 1558 7940
rect 1130 7760 1186 7816
rect 1254 7760 1310 7816
rect 1378 7760 1434 7816
rect 1502 7760 1558 7816
rect 1130 7636 1186 7692
rect 1254 7636 1310 7692
rect 1378 7636 1434 7692
rect 1502 7636 1558 7692
rect 85812 8008 85868 8064
rect 85936 8008 85992 8064
rect 86060 8008 86116 8064
rect 86184 8008 86240 8064
rect 85812 7884 85868 7940
rect 85936 7884 85992 7940
rect 86060 7884 86116 7940
rect 86184 7884 86240 7940
rect 85812 7760 85868 7816
rect 85936 7760 85992 7816
rect 86060 7760 86116 7816
rect 86184 7760 86240 7816
rect 85812 7636 85868 7692
rect 85936 7636 85992 7692
rect 86060 7636 86116 7692
rect 86184 7636 86240 7692
rect 86612 7108 86668 7164
rect 86736 7108 86792 7164
rect 86860 7108 86916 7164
rect 86984 7108 87040 7164
rect 1930 6984 1986 7040
rect 2054 6984 2110 7040
rect 2178 6984 2234 7040
rect 2302 6984 2358 7040
rect 1930 6860 1986 6916
rect 2054 6860 2110 6916
rect 2178 6860 2234 6916
rect 2302 6860 2358 6916
rect 86612 6984 86668 7040
rect 86736 6984 86792 7040
rect 86860 6984 86916 7040
rect 86984 6984 87040 7040
rect 86612 6860 86668 6916
rect 86736 6860 86792 6916
rect 86860 6860 86916 6916
rect 86984 6860 87040 6916
rect 86612 6736 86668 6792
rect 86736 6736 86792 6792
rect 86860 6736 86916 6792
rect 86984 6736 87040 6792
rect 1130 6208 1186 6264
rect 1254 6208 1310 6264
rect 1378 6208 1434 6264
rect 1502 6208 1558 6264
rect 1130 6084 1186 6140
rect 1254 6084 1310 6140
rect 1378 6084 1434 6140
rect 1502 6084 1558 6140
rect 1130 5960 1186 6016
rect 1254 5960 1310 6016
rect 1378 5960 1434 6016
rect 1502 5960 1558 6016
rect 1130 5836 1186 5892
rect 1254 5836 1310 5892
rect 1378 5836 1434 5892
rect 1502 5836 1558 5892
rect 85812 6208 85868 6264
rect 85936 6208 85992 6264
rect 86060 6208 86116 6264
rect 86184 6208 86240 6264
rect 85812 6084 85868 6140
rect 85936 6084 85992 6140
rect 86060 6084 86116 6140
rect 86184 6084 86240 6140
rect 85812 5960 85868 6016
rect 85936 5960 85992 6016
rect 86060 5960 86116 6016
rect 86184 5960 86240 6016
rect 85812 5836 85868 5892
rect 85936 5836 85992 5892
rect 86060 5836 86116 5892
rect 86184 5836 86240 5892
rect 86612 5308 86668 5364
rect 86736 5308 86792 5364
rect 86860 5308 86916 5364
rect 86984 5308 87040 5364
rect 1930 5184 1986 5240
rect 2054 5184 2110 5240
rect 2178 5184 2234 5240
rect 2302 5184 2358 5240
rect 1930 5060 1986 5116
rect 2054 5060 2110 5116
rect 2178 5060 2234 5116
rect 2302 5060 2358 5116
rect 86612 5184 86668 5240
rect 86736 5184 86792 5240
rect 86860 5184 86916 5240
rect 86984 5184 87040 5240
rect 86612 5060 86668 5116
rect 86736 5060 86792 5116
rect 86860 5060 86916 5116
rect 86984 5060 87040 5116
rect 86612 4936 86668 4992
rect 86736 4936 86792 4992
rect 86860 4936 86916 4992
rect 86984 4936 87040 4992
rect 1130 4408 1186 4464
rect 1254 4408 1310 4464
rect 1378 4408 1434 4464
rect 1502 4408 1558 4464
rect 1130 4284 1186 4340
rect 1254 4284 1310 4340
rect 1378 4284 1434 4340
rect 1502 4284 1558 4340
rect 1130 4160 1186 4216
rect 1254 4160 1310 4216
rect 1378 4160 1434 4216
rect 1502 4160 1558 4216
rect 1130 4036 1186 4092
rect 1254 4036 1310 4092
rect 1378 4036 1434 4092
rect 1502 4036 1558 4092
rect 85812 4408 85868 4464
rect 85936 4408 85992 4464
rect 86060 4408 86116 4464
rect 86184 4408 86240 4464
rect 85812 4284 85868 4340
rect 85936 4284 85992 4340
rect 86060 4284 86116 4340
rect 86184 4284 86240 4340
rect 85812 4160 85868 4216
rect 85936 4160 85992 4216
rect 86060 4160 86116 4216
rect 86184 4160 86240 4216
rect 85812 4036 85868 4092
rect 85936 4036 85992 4092
rect 86060 4036 86116 4092
rect 86184 4036 86240 4092
rect 86612 3576 86668 3632
rect 86736 3576 86792 3632
rect 86860 3576 86916 3632
rect 86984 3576 87040 3632
rect 1930 3384 1986 3440
rect 2054 3384 2110 3440
rect 2178 3384 2234 3440
rect 2302 3384 2358 3440
rect 1930 3260 1986 3316
rect 2054 3260 2110 3316
rect 2178 3260 2234 3316
rect 2302 3260 2358 3316
rect 86612 3452 86668 3508
rect 86736 3452 86792 3508
rect 86860 3452 86916 3508
rect 86984 3452 87040 3508
rect 86612 3328 86668 3384
rect 86736 3328 86792 3384
rect 86860 3328 86916 3384
rect 86984 3328 87040 3384
rect 86612 3204 86668 3260
rect 86736 3204 86792 3260
rect 86860 3204 86916 3260
rect 86984 3204 87040 3260
<< metal4 >>
rect 1044 85889 1644 95648
rect 1044 85833 1068 85889
rect 1124 85833 1192 85889
rect 1248 85833 1316 85889
rect 1372 85833 1440 85889
rect 1496 85833 1564 85889
rect 1620 85833 1644 85889
rect 1044 85765 1644 85833
rect 1044 85709 1068 85765
rect 1124 85709 1192 85765
rect 1248 85709 1316 85765
rect 1372 85709 1440 85765
rect 1496 85709 1564 85765
rect 1620 85709 1644 85765
rect 1044 85641 1644 85709
rect 1044 85585 1068 85641
rect 1124 85585 1192 85641
rect 1248 85585 1316 85641
rect 1372 85585 1440 85641
rect 1496 85585 1564 85641
rect 1620 85585 1644 85641
rect 1044 85517 1644 85585
rect 1044 85461 1068 85517
rect 1124 85461 1192 85517
rect 1248 85461 1316 85517
rect 1372 85461 1440 85517
rect 1496 85461 1564 85517
rect 1620 85461 1644 85517
rect 1044 85393 1644 85461
rect 1044 85337 1068 85393
rect 1124 85337 1192 85393
rect 1248 85337 1316 85393
rect 1372 85337 1440 85393
rect 1496 85337 1564 85393
rect 1620 85337 1644 85393
rect 1044 85269 1644 85337
rect 1044 85213 1068 85269
rect 1124 85213 1192 85269
rect 1248 85213 1316 85269
rect 1372 85213 1440 85269
rect 1496 85213 1564 85269
rect 1620 85213 1644 85269
rect 1044 85145 1644 85213
rect 1044 85089 1068 85145
rect 1124 85089 1192 85145
rect 1248 85089 1316 85145
rect 1372 85089 1440 85145
rect 1496 85089 1564 85145
rect 1620 85089 1644 85145
rect 1044 85021 1644 85089
rect 1044 84965 1068 85021
rect 1124 84965 1192 85021
rect 1248 84965 1316 85021
rect 1372 84965 1440 85021
rect 1496 84965 1564 85021
rect 1620 84965 1644 85021
rect 1044 84897 1644 84965
rect 1044 84841 1068 84897
rect 1124 84841 1192 84897
rect 1248 84841 1316 84897
rect 1372 84841 1440 84897
rect 1496 84841 1564 84897
rect 1620 84841 1644 84897
rect 1044 84773 1644 84841
rect 1044 84717 1068 84773
rect 1124 84717 1192 84773
rect 1248 84717 1316 84773
rect 1372 84717 1440 84773
rect 1496 84717 1564 84773
rect 1620 84717 1644 84773
rect 1044 84649 1644 84717
rect 1044 84593 1068 84649
rect 1124 84593 1192 84649
rect 1248 84593 1316 84649
rect 1372 84593 1440 84649
rect 1496 84593 1564 84649
rect 1620 84593 1644 84649
rect 1044 84525 1644 84593
rect 1044 84469 1068 84525
rect 1124 84469 1192 84525
rect 1248 84469 1316 84525
rect 1372 84469 1440 84525
rect 1496 84469 1564 84525
rect 1620 84469 1644 84525
rect 1044 84401 1644 84469
rect 1044 84345 1068 84401
rect 1124 84345 1192 84401
rect 1248 84345 1316 84401
rect 1372 84345 1440 84401
rect 1496 84345 1564 84401
rect 1620 84345 1644 84401
rect 1044 84277 1644 84345
rect 1044 84221 1068 84277
rect 1124 84221 1192 84277
rect 1248 84221 1316 84277
rect 1372 84221 1440 84277
rect 1496 84221 1564 84277
rect 1620 84221 1644 84277
rect 1044 84153 1644 84221
rect 1044 84097 1068 84153
rect 1124 84097 1192 84153
rect 1248 84097 1316 84153
rect 1372 84097 1440 84153
rect 1496 84097 1564 84153
rect 1620 84097 1644 84153
rect 1044 84029 1644 84097
rect 1044 83973 1068 84029
rect 1124 83973 1192 84029
rect 1248 83973 1316 84029
rect 1372 83973 1440 84029
rect 1496 83973 1564 84029
rect 1620 83973 1644 84029
rect 1044 83905 1644 83973
rect 1044 83849 1068 83905
rect 1124 83849 1192 83905
rect 1248 83849 1316 83905
rect 1372 83849 1440 83905
rect 1496 83849 1564 83905
rect 1620 83849 1644 83905
rect 1044 75000 1644 83849
rect 1044 74944 1068 75000
rect 1124 74944 1192 75000
rect 1248 74944 1316 75000
rect 1372 74944 1440 75000
rect 1496 74944 1564 75000
rect 1620 74944 1644 75000
rect 1044 74876 1644 74944
rect 1044 74820 1068 74876
rect 1124 74820 1192 74876
rect 1248 74820 1316 74876
rect 1372 74820 1440 74876
rect 1496 74820 1564 74876
rect 1620 74820 1644 74876
rect 1044 74752 1644 74820
rect 1044 74696 1068 74752
rect 1124 74696 1192 74752
rect 1248 74696 1316 74752
rect 1372 74696 1440 74752
rect 1496 74696 1564 74752
rect 1620 74696 1644 74752
rect 1044 74628 1644 74696
rect 1044 74572 1068 74628
rect 1124 74572 1192 74628
rect 1248 74572 1316 74628
rect 1372 74572 1440 74628
rect 1496 74572 1564 74628
rect 1620 74572 1644 74628
rect 1044 74504 1644 74572
rect 1044 74448 1068 74504
rect 1124 74448 1192 74504
rect 1248 74448 1316 74504
rect 1372 74448 1440 74504
rect 1496 74448 1564 74504
rect 1620 74448 1644 74504
rect 1044 74380 1644 74448
rect 1044 74324 1068 74380
rect 1124 74324 1192 74380
rect 1248 74324 1316 74380
rect 1372 74324 1440 74380
rect 1496 74324 1564 74380
rect 1620 74324 1644 74380
rect 1044 74256 1644 74324
rect 1044 74200 1068 74256
rect 1124 74200 1192 74256
rect 1248 74200 1316 74256
rect 1372 74200 1440 74256
rect 1496 74200 1564 74256
rect 1620 74200 1644 74256
rect 1044 74132 1644 74200
rect 1044 74076 1068 74132
rect 1124 74076 1192 74132
rect 1248 74076 1316 74132
rect 1372 74076 1440 74132
rect 1496 74076 1564 74132
rect 1620 74076 1644 74132
rect 1044 62064 1644 74076
rect 1044 62008 1130 62064
rect 1186 62008 1254 62064
rect 1310 62008 1378 62064
rect 1434 62008 1502 62064
rect 1558 62008 1644 62064
rect 1044 61940 1644 62008
rect 1044 61884 1130 61940
rect 1186 61884 1254 61940
rect 1310 61884 1378 61940
rect 1434 61884 1502 61940
rect 1558 61884 1644 61940
rect 1044 61816 1644 61884
rect 1044 61760 1130 61816
rect 1186 61760 1254 61816
rect 1310 61760 1378 61816
rect 1434 61760 1502 61816
rect 1558 61760 1644 61816
rect 1044 61692 1644 61760
rect 1044 61636 1130 61692
rect 1186 61636 1254 61692
rect 1310 61636 1378 61692
rect 1434 61636 1502 61692
rect 1558 61636 1644 61692
rect 1044 60264 1644 61636
rect 1044 60208 1130 60264
rect 1186 60208 1254 60264
rect 1310 60208 1378 60264
rect 1434 60208 1502 60264
rect 1558 60208 1644 60264
rect 1044 60140 1644 60208
rect 1044 60084 1130 60140
rect 1186 60084 1254 60140
rect 1310 60084 1378 60140
rect 1434 60084 1502 60140
rect 1558 60084 1644 60140
rect 1044 60016 1644 60084
rect 1044 59960 1130 60016
rect 1186 59960 1254 60016
rect 1310 59960 1378 60016
rect 1434 59960 1502 60016
rect 1558 59960 1644 60016
rect 1044 59892 1644 59960
rect 1044 59836 1130 59892
rect 1186 59836 1254 59892
rect 1310 59836 1378 59892
rect 1434 59836 1502 59892
rect 1558 59836 1644 59892
rect 1044 58464 1644 59836
rect 1044 58408 1130 58464
rect 1186 58408 1254 58464
rect 1310 58408 1378 58464
rect 1434 58408 1502 58464
rect 1558 58408 1644 58464
rect 1044 58340 1644 58408
rect 1044 58284 1130 58340
rect 1186 58284 1254 58340
rect 1310 58284 1378 58340
rect 1434 58284 1502 58340
rect 1558 58284 1644 58340
rect 1044 58216 1644 58284
rect 1044 58160 1130 58216
rect 1186 58160 1254 58216
rect 1310 58160 1378 58216
rect 1434 58160 1502 58216
rect 1558 58160 1644 58216
rect 1044 58092 1644 58160
rect 1044 58036 1130 58092
rect 1186 58036 1254 58092
rect 1310 58036 1378 58092
rect 1434 58036 1502 58092
rect 1558 58036 1644 58092
rect 1044 56664 1644 58036
rect 1044 56608 1130 56664
rect 1186 56608 1254 56664
rect 1310 56608 1378 56664
rect 1434 56608 1502 56664
rect 1558 56608 1644 56664
rect 1044 56540 1644 56608
rect 1044 56484 1130 56540
rect 1186 56484 1254 56540
rect 1310 56484 1378 56540
rect 1434 56484 1502 56540
rect 1558 56484 1644 56540
rect 1044 56416 1644 56484
rect 1044 56360 1130 56416
rect 1186 56360 1254 56416
rect 1310 56360 1378 56416
rect 1434 56360 1502 56416
rect 1558 56360 1644 56416
rect 1044 56292 1644 56360
rect 1044 56236 1130 56292
rect 1186 56236 1254 56292
rect 1310 56236 1378 56292
rect 1434 56236 1502 56292
rect 1558 56236 1644 56292
rect 1044 54864 1644 56236
rect 1044 54808 1130 54864
rect 1186 54808 1254 54864
rect 1310 54808 1378 54864
rect 1434 54808 1502 54864
rect 1558 54808 1644 54864
rect 1044 54740 1644 54808
rect 1044 54684 1130 54740
rect 1186 54684 1254 54740
rect 1310 54684 1378 54740
rect 1434 54684 1502 54740
rect 1558 54684 1644 54740
rect 1044 54616 1644 54684
rect 1044 54560 1130 54616
rect 1186 54560 1254 54616
rect 1310 54560 1378 54616
rect 1434 54560 1502 54616
rect 1558 54560 1644 54616
rect 1044 54492 1644 54560
rect 1044 54436 1130 54492
rect 1186 54436 1254 54492
rect 1310 54436 1378 54492
rect 1434 54436 1502 54492
rect 1558 54436 1644 54492
rect 1044 53064 1644 54436
rect 1044 53008 1130 53064
rect 1186 53008 1254 53064
rect 1310 53008 1378 53064
rect 1434 53008 1502 53064
rect 1558 53008 1644 53064
rect 1044 52940 1644 53008
rect 1044 52884 1130 52940
rect 1186 52884 1254 52940
rect 1310 52884 1378 52940
rect 1434 52884 1502 52940
rect 1558 52884 1644 52940
rect 1044 52816 1644 52884
rect 1044 52760 1130 52816
rect 1186 52760 1254 52816
rect 1310 52760 1378 52816
rect 1434 52760 1502 52816
rect 1558 52760 1644 52816
rect 1044 52692 1644 52760
rect 1044 52636 1130 52692
rect 1186 52636 1254 52692
rect 1310 52636 1378 52692
rect 1434 52636 1502 52692
rect 1558 52636 1644 52692
rect 1044 51264 1644 52636
rect 1044 51208 1130 51264
rect 1186 51208 1254 51264
rect 1310 51208 1378 51264
rect 1434 51208 1502 51264
rect 1558 51208 1644 51264
rect 1044 51140 1644 51208
rect 1044 51084 1130 51140
rect 1186 51084 1254 51140
rect 1310 51084 1378 51140
rect 1434 51084 1502 51140
rect 1558 51084 1644 51140
rect 1044 51016 1644 51084
rect 1044 50960 1130 51016
rect 1186 50960 1254 51016
rect 1310 50960 1378 51016
rect 1434 50960 1502 51016
rect 1558 50960 1644 51016
rect 1044 50892 1644 50960
rect 1044 50836 1130 50892
rect 1186 50836 1254 50892
rect 1310 50836 1378 50892
rect 1434 50836 1502 50892
rect 1558 50836 1644 50892
rect 1044 49464 1644 50836
rect 1044 49408 1130 49464
rect 1186 49408 1254 49464
rect 1310 49408 1378 49464
rect 1434 49408 1502 49464
rect 1558 49408 1644 49464
rect 1044 49340 1644 49408
rect 1044 49284 1130 49340
rect 1186 49284 1254 49340
rect 1310 49284 1378 49340
rect 1434 49284 1502 49340
rect 1558 49284 1644 49340
rect 1044 49216 1644 49284
rect 1044 49160 1130 49216
rect 1186 49160 1254 49216
rect 1310 49160 1378 49216
rect 1434 49160 1502 49216
rect 1558 49160 1644 49216
rect 1044 49092 1644 49160
rect 1044 49036 1130 49092
rect 1186 49036 1254 49092
rect 1310 49036 1378 49092
rect 1434 49036 1502 49092
rect 1558 49036 1644 49092
rect 1044 47664 1644 49036
rect 1044 47608 1130 47664
rect 1186 47608 1254 47664
rect 1310 47608 1378 47664
rect 1434 47608 1502 47664
rect 1558 47608 1644 47664
rect 1044 47540 1644 47608
rect 1044 47484 1130 47540
rect 1186 47484 1254 47540
rect 1310 47484 1378 47540
rect 1434 47484 1502 47540
rect 1558 47484 1644 47540
rect 1044 47416 1644 47484
rect 1044 47360 1130 47416
rect 1186 47360 1254 47416
rect 1310 47360 1378 47416
rect 1434 47360 1502 47416
rect 1558 47360 1644 47416
rect 1044 47292 1644 47360
rect 1044 47236 1130 47292
rect 1186 47236 1254 47292
rect 1310 47236 1378 47292
rect 1434 47236 1502 47292
rect 1558 47236 1644 47292
rect 1044 45864 1644 47236
rect 1044 45808 1130 45864
rect 1186 45808 1254 45864
rect 1310 45808 1378 45864
rect 1434 45808 1502 45864
rect 1558 45808 1644 45864
rect 1044 45740 1644 45808
rect 1044 45684 1130 45740
rect 1186 45684 1254 45740
rect 1310 45684 1378 45740
rect 1434 45684 1502 45740
rect 1558 45684 1644 45740
rect 1044 45616 1644 45684
rect 1044 45560 1130 45616
rect 1186 45560 1254 45616
rect 1310 45560 1378 45616
rect 1434 45560 1502 45616
rect 1558 45560 1644 45616
rect 1044 45492 1644 45560
rect 1044 45436 1130 45492
rect 1186 45436 1254 45492
rect 1310 45436 1378 45492
rect 1434 45436 1502 45492
rect 1558 45436 1644 45492
rect 1044 44064 1644 45436
rect 1044 44008 1130 44064
rect 1186 44008 1254 44064
rect 1310 44008 1378 44064
rect 1434 44008 1502 44064
rect 1558 44008 1644 44064
rect 1044 43940 1644 44008
rect 1044 43884 1130 43940
rect 1186 43884 1254 43940
rect 1310 43884 1378 43940
rect 1434 43884 1502 43940
rect 1558 43884 1644 43940
rect 1044 43816 1644 43884
rect 1044 43760 1130 43816
rect 1186 43760 1254 43816
rect 1310 43760 1378 43816
rect 1434 43760 1502 43816
rect 1558 43760 1644 43816
rect 1044 43692 1644 43760
rect 1044 43636 1130 43692
rect 1186 43636 1254 43692
rect 1310 43636 1378 43692
rect 1434 43636 1502 43692
rect 1558 43636 1644 43692
rect 1044 42264 1644 43636
rect 1044 42208 1130 42264
rect 1186 42208 1254 42264
rect 1310 42208 1378 42264
rect 1434 42208 1502 42264
rect 1558 42208 1644 42264
rect 1044 42140 1644 42208
rect 1044 42084 1130 42140
rect 1186 42084 1254 42140
rect 1310 42084 1378 42140
rect 1434 42084 1502 42140
rect 1558 42084 1644 42140
rect 1044 42016 1644 42084
rect 1044 41960 1130 42016
rect 1186 41960 1254 42016
rect 1310 41960 1378 42016
rect 1434 41960 1502 42016
rect 1558 41960 1644 42016
rect 1044 41892 1644 41960
rect 1044 41836 1130 41892
rect 1186 41836 1254 41892
rect 1310 41836 1378 41892
rect 1434 41836 1502 41892
rect 1558 41836 1644 41892
rect 1044 40464 1644 41836
rect 1044 40408 1130 40464
rect 1186 40408 1254 40464
rect 1310 40408 1378 40464
rect 1434 40408 1502 40464
rect 1558 40408 1644 40464
rect 1044 40340 1644 40408
rect 1044 40284 1130 40340
rect 1186 40284 1254 40340
rect 1310 40284 1378 40340
rect 1434 40284 1502 40340
rect 1558 40284 1644 40340
rect 1044 40216 1644 40284
rect 1044 40160 1130 40216
rect 1186 40160 1254 40216
rect 1310 40160 1378 40216
rect 1434 40160 1502 40216
rect 1558 40160 1644 40216
rect 1044 40092 1644 40160
rect 1044 40036 1130 40092
rect 1186 40036 1254 40092
rect 1310 40036 1378 40092
rect 1434 40036 1502 40092
rect 1558 40036 1644 40092
rect 1044 38664 1644 40036
rect 1044 38608 1130 38664
rect 1186 38608 1254 38664
rect 1310 38608 1378 38664
rect 1434 38608 1502 38664
rect 1558 38608 1644 38664
rect 1044 38540 1644 38608
rect 1044 38484 1130 38540
rect 1186 38484 1254 38540
rect 1310 38484 1378 38540
rect 1434 38484 1502 38540
rect 1558 38484 1644 38540
rect 1044 38416 1644 38484
rect 1044 38360 1130 38416
rect 1186 38360 1254 38416
rect 1310 38360 1378 38416
rect 1434 38360 1502 38416
rect 1558 38360 1644 38416
rect 1044 38292 1644 38360
rect 1044 38236 1130 38292
rect 1186 38236 1254 38292
rect 1310 38236 1378 38292
rect 1434 38236 1502 38292
rect 1558 38236 1644 38292
rect 1044 36864 1644 38236
rect 1044 36808 1130 36864
rect 1186 36808 1254 36864
rect 1310 36808 1378 36864
rect 1434 36808 1502 36864
rect 1558 36808 1644 36864
rect 1044 36740 1644 36808
rect 1044 36684 1130 36740
rect 1186 36684 1254 36740
rect 1310 36684 1378 36740
rect 1434 36684 1502 36740
rect 1558 36684 1644 36740
rect 1044 36616 1644 36684
rect 1044 36560 1130 36616
rect 1186 36560 1254 36616
rect 1310 36560 1378 36616
rect 1434 36560 1502 36616
rect 1558 36560 1644 36616
rect 1044 36492 1644 36560
rect 1044 36436 1130 36492
rect 1186 36436 1254 36492
rect 1310 36436 1378 36492
rect 1434 36436 1502 36492
rect 1558 36436 1644 36492
rect 1044 35064 1644 36436
rect 1044 35008 1130 35064
rect 1186 35008 1254 35064
rect 1310 35008 1378 35064
rect 1434 35008 1502 35064
rect 1558 35008 1644 35064
rect 1044 34940 1644 35008
rect 1044 34884 1130 34940
rect 1186 34884 1254 34940
rect 1310 34884 1378 34940
rect 1434 34884 1502 34940
rect 1558 34884 1644 34940
rect 1044 34816 1644 34884
rect 1044 34760 1130 34816
rect 1186 34760 1254 34816
rect 1310 34760 1378 34816
rect 1434 34760 1502 34816
rect 1558 34760 1644 34816
rect 1044 34692 1644 34760
rect 1044 34636 1130 34692
rect 1186 34636 1254 34692
rect 1310 34636 1378 34692
rect 1434 34636 1502 34692
rect 1558 34636 1644 34692
rect 1044 33264 1644 34636
rect 1044 33208 1130 33264
rect 1186 33208 1254 33264
rect 1310 33208 1378 33264
rect 1434 33208 1502 33264
rect 1558 33208 1644 33264
rect 1044 33140 1644 33208
rect 1044 33084 1130 33140
rect 1186 33084 1254 33140
rect 1310 33084 1378 33140
rect 1434 33084 1502 33140
rect 1558 33084 1644 33140
rect 1044 33016 1644 33084
rect 1044 32960 1130 33016
rect 1186 32960 1254 33016
rect 1310 32960 1378 33016
rect 1434 32960 1502 33016
rect 1558 32960 1644 33016
rect 1044 32892 1644 32960
rect 1044 32836 1130 32892
rect 1186 32836 1254 32892
rect 1310 32836 1378 32892
rect 1434 32836 1502 32892
rect 1558 32836 1644 32892
rect 1044 31464 1644 32836
rect 1044 31408 1130 31464
rect 1186 31408 1254 31464
rect 1310 31408 1378 31464
rect 1434 31408 1502 31464
rect 1558 31408 1644 31464
rect 1044 31340 1644 31408
rect 1044 31284 1130 31340
rect 1186 31284 1254 31340
rect 1310 31284 1378 31340
rect 1434 31284 1502 31340
rect 1558 31284 1644 31340
rect 1044 31216 1644 31284
rect 1044 31160 1130 31216
rect 1186 31160 1254 31216
rect 1310 31160 1378 31216
rect 1434 31160 1502 31216
rect 1558 31160 1644 31216
rect 1044 31092 1644 31160
rect 1044 31036 1130 31092
rect 1186 31036 1254 31092
rect 1310 31036 1378 31092
rect 1434 31036 1502 31092
rect 1558 31036 1644 31092
rect 1044 29664 1644 31036
rect 1044 29608 1130 29664
rect 1186 29608 1254 29664
rect 1310 29608 1378 29664
rect 1434 29608 1502 29664
rect 1558 29608 1644 29664
rect 1044 29540 1644 29608
rect 1044 29484 1130 29540
rect 1186 29484 1254 29540
rect 1310 29484 1378 29540
rect 1434 29484 1502 29540
rect 1558 29484 1644 29540
rect 1044 29416 1644 29484
rect 1044 29360 1130 29416
rect 1186 29360 1254 29416
rect 1310 29360 1378 29416
rect 1434 29360 1502 29416
rect 1558 29360 1644 29416
rect 1044 29292 1644 29360
rect 1044 29236 1130 29292
rect 1186 29236 1254 29292
rect 1310 29236 1378 29292
rect 1434 29236 1502 29292
rect 1558 29236 1644 29292
rect 1044 27864 1644 29236
rect 1044 27808 1130 27864
rect 1186 27808 1254 27864
rect 1310 27808 1378 27864
rect 1434 27808 1502 27864
rect 1558 27808 1644 27864
rect 1044 27740 1644 27808
rect 1044 27684 1130 27740
rect 1186 27684 1254 27740
rect 1310 27684 1378 27740
rect 1434 27684 1502 27740
rect 1558 27684 1644 27740
rect 1044 27616 1644 27684
rect 1044 27560 1130 27616
rect 1186 27560 1254 27616
rect 1310 27560 1378 27616
rect 1434 27560 1502 27616
rect 1558 27560 1644 27616
rect 1044 27492 1644 27560
rect 1044 27436 1130 27492
rect 1186 27436 1254 27492
rect 1310 27436 1378 27492
rect 1434 27436 1502 27492
rect 1558 27436 1644 27492
rect 1044 26064 1644 27436
rect 1044 26008 1130 26064
rect 1186 26008 1254 26064
rect 1310 26008 1378 26064
rect 1434 26008 1502 26064
rect 1558 26008 1644 26064
rect 1044 25940 1644 26008
rect 1044 25884 1130 25940
rect 1186 25884 1254 25940
rect 1310 25884 1378 25940
rect 1434 25884 1502 25940
rect 1558 25884 1644 25940
rect 1044 25816 1644 25884
rect 1044 25760 1130 25816
rect 1186 25760 1254 25816
rect 1310 25760 1378 25816
rect 1434 25760 1502 25816
rect 1558 25760 1644 25816
rect 1044 25692 1644 25760
rect 1044 25636 1130 25692
rect 1186 25636 1254 25692
rect 1310 25636 1378 25692
rect 1434 25636 1502 25692
rect 1558 25636 1644 25692
rect 1044 24264 1644 25636
rect 1044 24208 1130 24264
rect 1186 24208 1254 24264
rect 1310 24208 1378 24264
rect 1434 24208 1502 24264
rect 1558 24208 1644 24264
rect 1044 24140 1644 24208
rect 1044 24084 1130 24140
rect 1186 24084 1254 24140
rect 1310 24084 1378 24140
rect 1434 24084 1502 24140
rect 1558 24084 1644 24140
rect 1044 24016 1644 24084
rect 1044 23960 1130 24016
rect 1186 23960 1254 24016
rect 1310 23960 1378 24016
rect 1434 23960 1502 24016
rect 1558 23960 1644 24016
rect 1044 23892 1644 23960
rect 1044 23836 1130 23892
rect 1186 23836 1254 23892
rect 1310 23836 1378 23892
rect 1434 23836 1502 23892
rect 1558 23836 1644 23892
rect 1044 22464 1644 23836
rect 1044 22408 1130 22464
rect 1186 22408 1254 22464
rect 1310 22408 1378 22464
rect 1434 22408 1502 22464
rect 1558 22408 1644 22464
rect 1044 22340 1644 22408
rect 1044 22284 1130 22340
rect 1186 22284 1254 22340
rect 1310 22284 1378 22340
rect 1434 22284 1502 22340
rect 1558 22284 1644 22340
rect 1044 22216 1644 22284
rect 1044 22160 1130 22216
rect 1186 22160 1254 22216
rect 1310 22160 1378 22216
rect 1434 22160 1502 22216
rect 1558 22160 1644 22216
rect 1044 22092 1644 22160
rect 1044 22036 1130 22092
rect 1186 22036 1254 22092
rect 1310 22036 1378 22092
rect 1434 22036 1502 22092
rect 1558 22036 1644 22092
rect 1044 20664 1644 22036
rect 1044 20608 1130 20664
rect 1186 20608 1254 20664
rect 1310 20608 1378 20664
rect 1434 20608 1502 20664
rect 1558 20608 1644 20664
rect 1044 20540 1644 20608
rect 1044 20484 1130 20540
rect 1186 20484 1254 20540
rect 1310 20484 1378 20540
rect 1434 20484 1502 20540
rect 1558 20484 1644 20540
rect 1044 20416 1644 20484
rect 1044 20360 1130 20416
rect 1186 20360 1254 20416
rect 1310 20360 1378 20416
rect 1434 20360 1502 20416
rect 1558 20360 1644 20416
rect 1044 20292 1644 20360
rect 1044 20236 1130 20292
rect 1186 20236 1254 20292
rect 1310 20236 1378 20292
rect 1434 20236 1502 20292
rect 1558 20236 1644 20292
rect 1044 18864 1644 20236
rect 1044 18808 1130 18864
rect 1186 18808 1254 18864
rect 1310 18808 1378 18864
rect 1434 18808 1502 18864
rect 1558 18808 1644 18864
rect 1044 18740 1644 18808
rect 1044 18684 1130 18740
rect 1186 18684 1254 18740
rect 1310 18684 1378 18740
rect 1434 18684 1502 18740
rect 1558 18684 1644 18740
rect 1044 18616 1644 18684
rect 1044 18560 1130 18616
rect 1186 18560 1254 18616
rect 1310 18560 1378 18616
rect 1434 18560 1502 18616
rect 1558 18560 1644 18616
rect 1044 18492 1644 18560
rect 1044 18436 1130 18492
rect 1186 18436 1254 18492
rect 1310 18436 1378 18492
rect 1434 18436 1502 18492
rect 1558 18436 1644 18492
rect 1044 17064 1644 18436
rect 1044 17008 1130 17064
rect 1186 17008 1254 17064
rect 1310 17008 1378 17064
rect 1434 17008 1502 17064
rect 1558 17008 1644 17064
rect 1044 16940 1644 17008
rect 1044 16884 1130 16940
rect 1186 16884 1254 16940
rect 1310 16884 1378 16940
rect 1434 16884 1502 16940
rect 1558 16884 1644 16940
rect 1044 16816 1644 16884
rect 1044 16760 1130 16816
rect 1186 16760 1254 16816
rect 1310 16760 1378 16816
rect 1434 16760 1502 16816
rect 1558 16760 1644 16816
rect 1044 16692 1644 16760
rect 1044 16636 1130 16692
rect 1186 16636 1254 16692
rect 1310 16636 1378 16692
rect 1434 16636 1502 16692
rect 1558 16636 1644 16692
rect 1044 15264 1644 16636
rect 1044 15208 1130 15264
rect 1186 15208 1254 15264
rect 1310 15208 1378 15264
rect 1434 15208 1502 15264
rect 1558 15208 1644 15264
rect 1044 15140 1644 15208
rect 1044 15084 1130 15140
rect 1186 15084 1254 15140
rect 1310 15084 1378 15140
rect 1434 15084 1502 15140
rect 1558 15084 1644 15140
rect 1044 15016 1644 15084
rect 1044 14960 1130 15016
rect 1186 14960 1254 15016
rect 1310 14960 1378 15016
rect 1434 14960 1502 15016
rect 1558 14960 1644 15016
rect 1044 14892 1644 14960
rect 1044 14836 1130 14892
rect 1186 14836 1254 14892
rect 1310 14836 1378 14892
rect 1434 14836 1502 14892
rect 1558 14836 1644 14892
rect 1044 13464 1644 14836
rect 1044 13408 1130 13464
rect 1186 13408 1254 13464
rect 1310 13408 1378 13464
rect 1434 13408 1502 13464
rect 1558 13408 1644 13464
rect 1044 13340 1644 13408
rect 1044 13284 1130 13340
rect 1186 13284 1254 13340
rect 1310 13284 1378 13340
rect 1434 13284 1502 13340
rect 1558 13284 1644 13340
rect 1044 13216 1644 13284
rect 1044 13160 1130 13216
rect 1186 13160 1254 13216
rect 1310 13160 1378 13216
rect 1434 13160 1502 13216
rect 1558 13160 1644 13216
rect 1044 13092 1644 13160
rect 1044 13036 1130 13092
rect 1186 13036 1254 13092
rect 1310 13036 1378 13092
rect 1434 13036 1502 13092
rect 1558 13036 1644 13092
rect 1044 11664 1644 13036
rect 1044 11608 1130 11664
rect 1186 11608 1254 11664
rect 1310 11608 1378 11664
rect 1434 11608 1502 11664
rect 1558 11608 1644 11664
rect 1044 11540 1644 11608
rect 1044 11484 1130 11540
rect 1186 11484 1254 11540
rect 1310 11484 1378 11540
rect 1434 11484 1502 11540
rect 1558 11484 1644 11540
rect 1044 11416 1644 11484
rect 1044 11360 1130 11416
rect 1186 11360 1254 11416
rect 1310 11360 1378 11416
rect 1434 11360 1502 11416
rect 1558 11360 1644 11416
rect 1044 11292 1644 11360
rect 1044 11236 1130 11292
rect 1186 11236 1254 11292
rect 1310 11236 1378 11292
rect 1434 11236 1502 11292
rect 1558 11236 1644 11292
rect 1044 9864 1644 11236
rect 1044 9808 1130 9864
rect 1186 9808 1254 9864
rect 1310 9808 1378 9864
rect 1434 9808 1502 9864
rect 1558 9808 1644 9864
rect 1044 9740 1644 9808
rect 1044 9684 1130 9740
rect 1186 9684 1254 9740
rect 1310 9684 1378 9740
rect 1434 9684 1502 9740
rect 1558 9684 1644 9740
rect 1044 9616 1644 9684
rect 1044 9560 1130 9616
rect 1186 9560 1254 9616
rect 1310 9560 1378 9616
rect 1434 9560 1502 9616
rect 1558 9560 1644 9616
rect 1044 9492 1644 9560
rect 1044 9436 1130 9492
rect 1186 9436 1254 9492
rect 1310 9436 1378 9492
rect 1434 9436 1502 9492
rect 1558 9436 1644 9492
rect 1044 8064 1644 9436
rect 1044 8008 1130 8064
rect 1186 8008 1254 8064
rect 1310 8008 1378 8064
rect 1434 8008 1502 8064
rect 1558 8008 1644 8064
rect 1044 7940 1644 8008
rect 1044 7884 1130 7940
rect 1186 7884 1254 7940
rect 1310 7884 1378 7940
rect 1434 7884 1502 7940
rect 1558 7884 1644 7940
rect 1044 7816 1644 7884
rect 1044 7760 1130 7816
rect 1186 7760 1254 7816
rect 1310 7760 1378 7816
rect 1434 7760 1502 7816
rect 1558 7760 1644 7816
rect 1044 7692 1644 7760
rect 1044 7636 1130 7692
rect 1186 7636 1254 7692
rect 1310 7636 1378 7692
rect 1434 7636 1502 7692
rect 1558 7636 1644 7692
rect 1044 6264 1644 7636
rect 1044 6208 1130 6264
rect 1186 6208 1254 6264
rect 1310 6208 1378 6264
rect 1434 6208 1502 6264
rect 1558 6208 1644 6264
rect 1044 6140 1644 6208
rect 1044 6084 1130 6140
rect 1186 6084 1254 6140
rect 1310 6084 1378 6140
rect 1434 6084 1502 6140
rect 1558 6084 1644 6140
rect 1044 6016 1644 6084
rect 1044 5960 1130 6016
rect 1186 5960 1254 6016
rect 1310 5960 1378 6016
rect 1434 5960 1502 6016
rect 1558 5960 1644 6016
rect 1044 5892 1644 5960
rect 1044 5836 1130 5892
rect 1186 5836 1254 5892
rect 1310 5836 1378 5892
rect 1434 5836 1502 5892
rect 1558 5836 1644 5892
rect 1044 4464 1644 5836
rect 1044 4408 1130 4464
rect 1186 4408 1254 4464
rect 1310 4408 1378 4464
rect 1434 4408 1502 4464
rect 1558 4408 1644 4464
rect 1044 4340 1644 4408
rect 1044 4284 1130 4340
rect 1186 4284 1254 4340
rect 1310 4284 1378 4340
rect 1434 4284 1502 4340
rect 1558 4284 1644 4340
rect 1044 4216 1644 4284
rect 1044 4160 1130 4216
rect 1186 4160 1254 4216
rect 1310 4160 1378 4216
rect 1434 4160 1502 4216
rect 1558 4160 1644 4216
rect 1044 4092 1644 4160
rect 1044 4036 1130 4092
rect 1186 4036 1254 4092
rect 1310 4036 1378 4092
rect 1434 4036 1502 4092
rect 1558 4036 1644 4092
rect 1044 3136 1644 4036
rect 1844 95425 2444 95648
rect 1844 95369 1901 95425
rect 1957 95369 2444 95425
rect 1844 95301 2444 95369
rect 1844 95245 1901 95301
rect 1957 95245 2444 95301
rect 1844 95177 2444 95245
rect 1844 95121 1901 95177
rect 1957 95121 2444 95177
rect 1844 95053 2444 95121
rect 1844 94997 1901 95053
rect 1957 94997 2444 95053
rect 1844 94929 2444 94997
rect 1844 94873 1901 94929
rect 1957 94873 2444 94929
rect 1844 94805 2444 94873
rect 1844 94749 1901 94805
rect 1957 94749 2444 94805
rect 1844 94681 2444 94749
rect 1844 94625 1901 94681
rect 1957 94625 2444 94681
rect 1844 94557 2444 94625
rect 1844 94501 1901 94557
rect 1957 94501 2444 94557
rect 1844 94433 2444 94501
rect 1844 94377 1901 94433
rect 1957 94377 2444 94433
rect 1844 94309 2444 94377
rect 1844 94253 1901 94309
rect 1957 94253 2444 94309
rect 1844 90901 2444 94253
rect 1844 90845 1930 90901
rect 1986 90845 2054 90901
rect 2110 90845 2178 90901
rect 2234 90845 2302 90901
rect 2358 90845 2444 90901
rect 1844 90777 2444 90845
rect 1844 90721 1930 90777
rect 1986 90721 2054 90777
rect 2110 90721 2178 90777
rect 2234 90721 2302 90777
rect 2358 90721 2444 90777
rect 1844 90653 2444 90721
rect 1844 90597 1930 90653
rect 1986 90597 2054 90653
rect 2110 90597 2178 90653
rect 2234 90597 2302 90653
rect 2358 90597 2444 90653
rect 1844 90529 2444 90597
rect 1844 90473 1930 90529
rect 1986 90473 2054 90529
rect 2110 90473 2178 90529
rect 2234 90473 2302 90529
rect 2358 90473 2444 90529
rect 1844 83587 2444 90473
rect 1844 83531 1868 83587
rect 1924 83531 1992 83587
rect 2048 83531 2116 83587
rect 2172 83531 2240 83587
rect 2296 83531 2364 83587
rect 2420 83531 2444 83587
rect 1844 83463 2444 83531
rect 1844 83407 1868 83463
rect 1924 83407 1992 83463
rect 2048 83407 2116 83463
rect 2172 83407 2240 83463
rect 2296 83407 2364 83463
rect 2420 83407 2444 83463
rect 1844 83339 2444 83407
rect 1844 83283 1868 83339
rect 1924 83283 1992 83339
rect 2048 83283 2116 83339
rect 2172 83283 2240 83339
rect 2296 83283 2364 83339
rect 2420 83283 2444 83339
rect 1844 83215 2444 83283
rect 1844 83159 1868 83215
rect 1924 83159 1992 83215
rect 2048 83159 2116 83215
rect 2172 83159 2240 83215
rect 2296 83159 2364 83215
rect 2420 83159 2444 83215
rect 1844 83091 2444 83159
rect 1844 83035 1868 83091
rect 1924 83035 1992 83091
rect 2048 83035 2116 83091
rect 2172 83035 2240 83091
rect 2296 83035 2364 83091
rect 2420 83035 2444 83091
rect 1844 82967 2444 83035
rect 1844 82911 1868 82967
rect 1924 82911 1992 82967
rect 2048 82911 2116 82967
rect 2172 82911 2240 82967
rect 2296 82911 2364 82967
rect 2420 82911 2444 82967
rect 1844 82843 2444 82911
rect 1844 82787 1868 82843
rect 1924 82787 1992 82843
rect 2048 82787 2116 82843
rect 2172 82787 2240 82843
rect 2296 82787 2364 82843
rect 2420 82787 2444 82843
rect 1844 82719 2444 82787
rect 1844 82663 1868 82719
rect 1924 82663 1992 82719
rect 2048 82663 2116 82719
rect 2172 82663 2240 82719
rect 2296 82663 2364 82719
rect 2420 82663 2444 82719
rect 1844 82595 2444 82663
rect 1844 82539 1868 82595
rect 1924 82539 1992 82595
rect 2048 82539 2116 82595
rect 2172 82539 2240 82595
rect 2296 82539 2364 82595
rect 2420 82539 2444 82595
rect 1844 82471 2444 82539
rect 1844 82415 1868 82471
rect 1924 82415 1992 82471
rect 2048 82415 2116 82471
rect 2172 82415 2240 82471
rect 2296 82415 2364 82471
rect 2420 82415 2444 82471
rect 1844 82347 2444 82415
rect 1844 82291 1868 82347
rect 1924 82291 1992 82347
rect 2048 82291 2116 82347
rect 2172 82291 2240 82347
rect 2296 82291 2364 82347
rect 2420 82291 2444 82347
rect 1844 82223 2444 82291
rect 1844 82167 1868 82223
rect 1924 82167 1992 82223
rect 2048 82167 2116 82223
rect 2172 82167 2240 82223
rect 2296 82167 2364 82223
rect 2420 82167 2444 82223
rect 1844 82099 2444 82167
rect 1844 82043 1868 82099
rect 1924 82043 1992 82099
rect 2048 82043 2116 82099
rect 2172 82043 2240 82099
rect 2296 82043 2364 82099
rect 2420 82043 2444 82099
rect 1844 81975 2444 82043
rect 1844 81919 1868 81975
rect 1924 81919 1992 81975
rect 2048 81919 2116 81975
rect 2172 81919 2240 81975
rect 2296 81919 2364 81975
rect 2420 81919 2444 81975
rect 1844 81851 2444 81919
rect 1844 81795 1868 81851
rect 1924 81795 1992 81851
rect 2048 81795 2116 81851
rect 2172 81795 2240 81851
rect 2296 81795 2364 81851
rect 2420 81795 2444 81851
rect 1844 81727 2444 81795
rect 1844 81671 1868 81727
rect 1924 81671 1992 81727
rect 2048 81671 2116 81727
rect 2172 81671 2240 81727
rect 2296 81671 2364 81727
rect 2420 81671 2444 81727
rect 1844 81603 2444 81671
rect 1844 81547 1868 81603
rect 1924 81547 1992 81603
rect 2048 81547 2116 81603
rect 2172 81547 2240 81603
rect 2296 81547 2364 81603
rect 2420 81547 2444 81603
rect 1844 81479 2444 81547
rect 1844 81423 1868 81479
rect 1924 81423 1992 81479
rect 2048 81423 2116 81479
rect 2172 81423 2240 81479
rect 2296 81423 2364 81479
rect 2420 81423 2444 81479
rect 1844 81355 2444 81423
rect 1844 81299 1868 81355
rect 1924 81299 1992 81355
rect 2048 81299 2116 81355
rect 2172 81299 2240 81355
rect 2296 81299 2364 81355
rect 2420 81299 2444 81355
rect 1844 81231 2444 81299
rect 1844 81175 1868 81231
rect 1924 81175 1992 81231
rect 2048 81175 2116 81231
rect 2172 81175 2240 81231
rect 2296 81175 2364 81231
rect 2420 81175 2444 81231
rect 1844 81107 2444 81175
rect 1844 81051 1868 81107
rect 1924 81051 1992 81107
rect 2048 81051 2116 81107
rect 2172 81051 2240 81107
rect 2296 81051 2364 81107
rect 2420 81051 2444 81107
rect 1844 80983 2444 81051
rect 1844 80927 1868 80983
rect 1924 80927 1992 80983
rect 2048 80927 2116 80983
rect 2172 80927 2240 80983
rect 2296 80927 2364 80983
rect 2420 80927 2444 80983
rect 1844 80859 2444 80927
rect 1844 80803 1868 80859
rect 1924 80803 1992 80859
rect 2048 80803 2116 80859
rect 2172 80803 2240 80859
rect 2296 80803 2364 80859
rect 2420 80803 2444 80859
rect 1844 80735 2444 80803
rect 1844 80679 1868 80735
rect 1924 80679 1992 80735
rect 2048 80679 2116 80735
rect 2172 80679 2240 80735
rect 2296 80679 2364 80735
rect 2420 80679 2444 80735
rect 1844 80611 2444 80679
rect 1844 80555 1868 80611
rect 1924 80555 1992 80611
rect 2048 80555 2116 80611
rect 2172 80555 2240 80611
rect 2296 80555 2364 80611
rect 2420 80555 2444 80611
rect 1844 80487 2444 80555
rect 1844 80431 1868 80487
rect 1924 80431 1992 80487
rect 2048 80431 2116 80487
rect 2172 80431 2240 80487
rect 2296 80431 2364 80487
rect 2420 80431 2444 80487
rect 1844 80363 2444 80431
rect 1844 80307 1868 80363
rect 1924 80307 1992 80363
rect 2048 80307 2116 80363
rect 2172 80307 2240 80363
rect 2296 80307 2364 80363
rect 2420 80307 2444 80363
rect 1844 63414 2444 80307
rect 1844 63358 1930 63414
rect 1986 63358 2054 63414
rect 2110 63358 2178 63414
rect 2234 63358 2302 63414
rect 2358 63358 2444 63414
rect 1844 63290 2444 63358
rect 1844 63234 1930 63290
rect 1986 63234 2054 63290
rect 2110 63234 2178 63290
rect 2234 63234 2302 63290
rect 2358 63234 2444 63290
rect 1844 63166 2444 63234
rect 1844 63110 1930 63166
rect 1986 63110 2054 63166
rect 2110 63110 2178 63166
rect 2234 63110 2302 63166
rect 2358 63110 2444 63166
rect 1844 63042 2444 63110
rect 1844 62986 1930 63042
rect 1986 62986 2054 63042
rect 2110 62986 2178 63042
rect 2234 62986 2302 63042
rect 2358 62986 2444 63042
rect 1844 62840 2444 62986
rect 1844 62784 1930 62840
rect 1986 62784 2054 62840
rect 2110 62784 2178 62840
rect 2234 62784 2302 62840
rect 2358 62784 2444 62840
rect 1844 62716 2444 62784
rect 1844 62660 1930 62716
rect 1986 62660 2054 62716
rect 2110 62660 2178 62716
rect 2234 62660 2302 62716
rect 2358 62660 2444 62716
rect 1844 61040 2444 62660
rect 1844 60984 1930 61040
rect 1986 60984 2054 61040
rect 2110 60984 2178 61040
rect 2234 60984 2302 61040
rect 2358 60984 2444 61040
rect 1844 60916 2444 60984
rect 1844 60860 1930 60916
rect 1986 60860 2054 60916
rect 2110 60860 2178 60916
rect 2234 60860 2302 60916
rect 2358 60860 2444 60916
rect 1844 59240 2444 60860
rect 1844 59184 1930 59240
rect 1986 59184 2054 59240
rect 2110 59184 2178 59240
rect 2234 59184 2302 59240
rect 2358 59184 2444 59240
rect 1844 59116 2444 59184
rect 1844 59060 1930 59116
rect 1986 59060 2054 59116
rect 2110 59060 2178 59116
rect 2234 59060 2302 59116
rect 2358 59060 2444 59116
rect 1844 57440 2444 59060
rect 1844 57384 1930 57440
rect 1986 57384 2054 57440
rect 2110 57384 2178 57440
rect 2234 57384 2302 57440
rect 2358 57384 2444 57440
rect 1844 57316 2444 57384
rect 1844 57260 1930 57316
rect 1986 57260 2054 57316
rect 2110 57260 2178 57316
rect 2234 57260 2302 57316
rect 2358 57260 2444 57316
rect 1844 55640 2444 57260
rect 1844 55584 1930 55640
rect 1986 55584 2054 55640
rect 2110 55584 2178 55640
rect 2234 55584 2302 55640
rect 2358 55584 2444 55640
rect 1844 55516 2444 55584
rect 1844 55460 1930 55516
rect 1986 55460 2054 55516
rect 2110 55460 2178 55516
rect 2234 55460 2302 55516
rect 2358 55460 2444 55516
rect 1844 53840 2444 55460
rect 1844 53784 1930 53840
rect 1986 53784 2054 53840
rect 2110 53784 2178 53840
rect 2234 53784 2302 53840
rect 2358 53784 2444 53840
rect 1844 53716 2444 53784
rect 1844 53660 1930 53716
rect 1986 53660 2054 53716
rect 2110 53660 2178 53716
rect 2234 53660 2302 53716
rect 2358 53660 2444 53716
rect 1844 52040 2444 53660
rect 1844 51984 1930 52040
rect 1986 51984 2054 52040
rect 2110 51984 2178 52040
rect 2234 51984 2302 52040
rect 2358 51984 2444 52040
rect 1844 51916 2444 51984
rect 1844 51860 1930 51916
rect 1986 51860 2054 51916
rect 2110 51860 2178 51916
rect 2234 51860 2302 51916
rect 2358 51860 2444 51916
rect 1844 50240 2444 51860
rect 1844 50184 1930 50240
rect 1986 50184 2054 50240
rect 2110 50184 2178 50240
rect 2234 50184 2302 50240
rect 2358 50184 2444 50240
rect 1844 50116 2444 50184
rect 1844 50060 1930 50116
rect 1986 50060 2054 50116
rect 2110 50060 2178 50116
rect 2234 50060 2302 50116
rect 2358 50060 2444 50116
rect 1844 48440 2444 50060
rect 1844 48384 1930 48440
rect 1986 48384 2054 48440
rect 2110 48384 2178 48440
rect 2234 48384 2302 48440
rect 2358 48384 2444 48440
rect 1844 48316 2444 48384
rect 1844 48260 1930 48316
rect 1986 48260 2054 48316
rect 2110 48260 2178 48316
rect 2234 48260 2302 48316
rect 2358 48260 2444 48316
rect 1844 46640 2444 48260
rect 1844 46584 1930 46640
rect 1986 46584 2054 46640
rect 2110 46584 2178 46640
rect 2234 46584 2302 46640
rect 2358 46584 2444 46640
rect 1844 46516 2444 46584
rect 1844 46460 1930 46516
rect 1986 46460 2054 46516
rect 2110 46460 2178 46516
rect 2234 46460 2302 46516
rect 2358 46460 2444 46516
rect 1844 44840 2444 46460
rect 1844 44784 1930 44840
rect 1986 44784 2054 44840
rect 2110 44784 2178 44840
rect 2234 44784 2302 44840
rect 2358 44784 2444 44840
rect 1844 44716 2444 44784
rect 1844 44660 1930 44716
rect 1986 44660 2054 44716
rect 2110 44660 2178 44716
rect 2234 44660 2302 44716
rect 2358 44660 2444 44716
rect 1844 43040 2444 44660
rect 1844 42984 1930 43040
rect 1986 42984 2054 43040
rect 2110 42984 2178 43040
rect 2234 42984 2302 43040
rect 2358 42984 2444 43040
rect 1844 42916 2444 42984
rect 1844 42860 1930 42916
rect 1986 42860 2054 42916
rect 2110 42860 2178 42916
rect 2234 42860 2302 42916
rect 2358 42860 2444 42916
rect 1844 41240 2444 42860
rect 1844 41184 1930 41240
rect 1986 41184 2054 41240
rect 2110 41184 2178 41240
rect 2234 41184 2302 41240
rect 2358 41184 2444 41240
rect 1844 41116 2444 41184
rect 1844 41060 1930 41116
rect 1986 41060 2054 41116
rect 2110 41060 2178 41116
rect 2234 41060 2302 41116
rect 2358 41060 2444 41116
rect 1844 39440 2444 41060
rect 1844 39384 1930 39440
rect 1986 39384 2054 39440
rect 2110 39384 2178 39440
rect 2234 39384 2302 39440
rect 2358 39384 2444 39440
rect 1844 39316 2444 39384
rect 1844 39260 1930 39316
rect 1986 39260 2054 39316
rect 2110 39260 2178 39316
rect 2234 39260 2302 39316
rect 2358 39260 2444 39316
rect 1844 37640 2444 39260
rect 1844 37584 1930 37640
rect 1986 37584 2054 37640
rect 2110 37584 2178 37640
rect 2234 37584 2302 37640
rect 2358 37584 2444 37640
rect 1844 37516 2444 37584
rect 1844 37460 1930 37516
rect 1986 37460 2054 37516
rect 2110 37460 2178 37516
rect 2234 37460 2302 37516
rect 2358 37460 2444 37516
rect 1844 35840 2444 37460
rect 1844 35784 1930 35840
rect 1986 35784 2054 35840
rect 2110 35784 2178 35840
rect 2234 35784 2302 35840
rect 2358 35784 2444 35840
rect 1844 35716 2444 35784
rect 1844 35660 1930 35716
rect 1986 35660 2054 35716
rect 2110 35660 2178 35716
rect 2234 35660 2302 35716
rect 2358 35660 2444 35716
rect 1844 34040 2444 35660
rect 1844 33984 1930 34040
rect 1986 33984 2054 34040
rect 2110 33984 2178 34040
rect 2234 33984 2302 34040
rect 2358 33984 2444 34040
rect 1844 33916 2444 33984
rect 1844 33860 1930 33916
rect 1986 33860 2054 33916
rect 2110 33860 2178 33916
rect 2234 33860 2302 33916
rect 2358 33860 2444 33916
rect 1844 32240 2444 33860
rect 1844 32184 1930 32240
rect 1986 32184 2054 32240
rect 2110 32184 2178 32240
rect 2234 32184 2302 32240
rect 2358 32184 2444 32240
rect 1844 32116 2444 32184
rect 1844 32060 1930 32116
rect 1986 32060 2054 32116
rect 2110 32060 2178 32116
rect 2234 32060 2302 32116
rect 2358 32060 2444 32116
rect 1844 30440 2444 32060
rect 1844 30384 1930 30440
rect 1986 30384 2054 30440
rect 2110 30384 2178 30440
rect 2234 30384 2302 30440
rect 2358 30384 2444 30440
rect 1844 30316 2444 30384
rect 1844 30260 1930 30316
rect 1986 30260 2054 30316
rect 2110 30260 2178 30316
rect 2234 30260 2302 30316
rect 2358 30260 2444 30316
rect 1844 28640 2444 30260
rect 1844 28584 1930 28640
rect 1986 28584 2054 28640
rect 2110 28584 2178 28640
rect 2234 28584 2302 28640
rect 2358 28584 2444 28640
rect 1844 28516 2444 28584
rect 1844 28460 1930 28516
rect 1986 28460 2054 28516
rect 2110 28460 2178 28516
rect 2234 28460 2302 28516
rect 2358 28460 2444 28516
rect 1844 26840 2444 28460
rect 1844 26784 1930 26840
rect 1986 26784 2054 26840
rect 2110 26784 2178 26840
rect 2234 26784 2302 26840
rect 2358 26784 2444 26840
rect 1844 26716 2444 26784
rect 1844 26660 1930 26716
rect 1986 26660 2054 26716
rect 2110 26660 2178 26716
rect 2234 26660 2302 26716
rect 2358 26660 2444 26716
rect 1844 25040 2444 26660
rect 1844 24984 1930 25040
rect 1986 24984 2054 25040
rect 2110 24984 2178 25040
rect 2234 24984 2302 25040
rect 2358 24984 2444 25040
rect 1844 24916 2444 24984
rect 1844 24860 1930 24916
rect 1986 24860 2054 24916
rect 2110 24860 2178 24916
rect 2234 24860 2302 24916
rect 2358 24860 2444 24916
rect 1844 23240 2444 24860
rect 1844 23184 1930 23240
rect 1986 23184 2054 23240
rect 2110 23184 2178 23240
rect 2234 23184 2302 23240
rect 2358 23184 2444 23240
rect 1844 23116 2444 23184
rect 1844 23060 1930 23116
rect 1986 23060 2054 23116
rect 2110 23060 2178 23116
rect 2234 23060 2302 23116
rect 2358 23060 2444 23116
rect 1844 21440 2444 23060
rect 1844 21384 1930 21440
rect 1986 21384 2054 21440
rect 2110 21384 2178 21440
rect 2234 21384 2302 21440
rect 2358 21384 2444 21440
rect 1844 21316 2444 21384
rect 1844 21260 1930 21316
rect 1986 21260 2054 21316
rect 2110 21260 2178 21316
rect 2234 21260 2302 21316
rect 2358 21260 2444 21316
rect 1844 19640 2444 21260
rect 1844 19584 1930 19640
rect 1986 19584 2054 19640
rect 2110 19584 2178 19640
rect 2234 19584 2302 19640
rect 2358 19584 2444 19640
rect 1844 19516 2444 19584
rect 1844 19460 1930 19516
rect 1986 19460 2054 19516
rect 2110 19460 2178 19516
rect 2234 19460 2302 19516
rect 2358 19460 2444 19516
rect 1844 17840 2444 19460
rect 1844 17784 1930 17840
rect 1986 17784 2054 17840
rect 2110 17784 2178 17840
rect 2234 17784 2302 17840
rect 2358 17784 2444 17840
rect 1844 17716 2444 17784
rect 1844 17660 1930 17716
rect 1986 17660 2054 17716
rect 2110 17660 2178 17716
rect 2234 17660 2302 17716
rect 2358 17660 2444 17716
rect 1844 16040 2444 17660
rect 1844 15984 1930 16040
rect 1986 15984 2054 16040
rect 2110 15984 2178 16040
rect 2234 15984 2302 16040
rect 2358 15984 2444 16040
rect 1844 15916 2444 15984
rect 1844 15860 1930 15916
rect 1986 15860 2054 15916
rect 2110 15860 2178 15916
rect 2234 15860 2302 15916
rect 2358 15860 2444 15916
rect 1844 14240 2444 15860
rect 1844 14184 1930 14240
rect 1986 14184 2054 14240
rect 2110 14184 2178 14240
rect 2234 14184 2302 14240
rect 2358 14184 2444 14240
rect 1844 14116 2444 14184
rect 1844 14060 1930 14116
rect 1986 14060 2054 14116
rect 2110 14060 2178 14116
rect 2234 14060 2302 14116
rect 2358 14060 2444 14116
rect 1844 12440 2444 14060
rect 1844 12384 1930 12440
rect 1986 12384 2054 12440
rect 2110 12384 2178 12440
rect 2234 12384 2302 12440
rect 2358 12384 2444 12440
rect 1844 12316 2444 12384
rect 1844 12260 1930 12316
rect 1986 12260 2054 12316
rect 2110 12260 2178 12316
rect 2234 12260 2302 12316
rect 2358 12260 2444 12316
rect 1844 10640 2444 12260
rect 1844 10584 1930 10640
rect 1986 10584 2054 10640
rect 2110 10584 2178 10640
rect 2234 10584 2302 10640
rect 2358 10584 2444 10640
rect 1844 10516 2444 10584
rect 1844 10460 1930 10516
rect 1986 10460 2054 10516
rect 2110 10460 2178 10516
rect 2234 10460 2302 10516
rect 2358 10460 2444 10516
rect 1844 8840 2444 10460
rect 1844 8784 1930 8840
rect 1986 8784 2054 8840
rect 2110 8784 2178 8840
rect 2234 8784 2302 8840
rect 2358 8784 2444 8840
rect 1844 8716 2444 8784
rect 1844 8660 1930 8716
rect 1986 8660 2054 8716
rect 2110 8660 2178 8716
rect 2234 8660 2302 8716
rect 2358 8660 2444 8716
rect 1844 7040 2444 8660
rect 1844 6984 1930 7040
rect 1986 6984 2054 7040
rect 2110 6984 2178 7040
rect 2234 6984 2302 7040
rect 2358 6984 2444 7040
rect 1844 6916 2444 6984
rect 1844 6860 1930 6916
rect 1986 6860 2054 6916
rect 2110 6860 2178 6916
rect 2234 6860 2302 6916
rect 2358 6860 2444 6916
rect 1844 5240 2444 6860
rect 1844 5184 1930 5240
rect 1986 5184 2054 5240
rect 2110 5184 2178 5240
rect 2234 5184 2302 5240
rect 2358 5184 2444 5240
rect 1844 5116 2444 5184
rect 1844 5060 1930 5116
rect 1986 5060 2054 5116
rect 2110 5060 2178 5116
rect 2234 5060 2302 5116
rect 2358 5060 2444 5116
rect 1844 3440 2444 5060
rect 1844 3384 1930 3440
rect 1986 3384 2054 3440
rect 2110 3384 2178 3440
rect 2234 3384 2302 3440
rect 2358 3384 2444 3440
rect 1844 3316 2444 3384
rect 1844 3260 1930 3316
rect 1986 3260 2054 3316
rect 2110 3260 2178 3316
rect 2234 3260 2302 3316
rect 2358 3260 2444 3316
rect 1844 3136 2444 3260
rect 85726 89791 86326 95648
rect 85726 89735 85750 89791
rect 85806 89735 85874 89791
rect 85930 89735 85998 89791
rect 86054 89735 86122 89791
rect 86178 89735 86246 89791
rect 86302 89735 86326 89791
rect 85726 89667 86326 89735
rect 85726 89611 85750 89667
rect 85806 89611 85874 89667
rect 85930 89611 85998 89667
rect 86054 89611 86122 89667
rect 86178 89611 86246 89667
rect 86302 89611 86326 89667
rect 85726 89543 86326 89611
rect 85726 89487 85750 89543
rect 85806 89487 85874 89543
rect 85930 89487 85998 89543
rect 86054 89487 86122 89543
rect 86178 89487 86246 89543
rect 86302 89487 86326 89543
rect 85726 89419 86326 89487
rect 85726 89363 85750 89419
rect 85806 89363 85874 89419
rect 85930 89363 85998 89419
rect 86054 89363 86122 89419
rect 86178 89363 86246 89419
rect 86302 89363 86326 89419
rect 85726 89295 86326 89363
rect 85726 89239 85750 89295
rect 85806 89239 85874 89295
rect 85930 89239 85998 89295
rect 86054 89239 86122 89295
rect 86178 89239 86246 89295
rect 86302 89239 86326 89295
rect 85726 89171 86326 89239
rect 85726 89115 85750 89171
rect 85806 89115 85874 89171
rect 85930 89115 85998 89171
rect 86054 89115 86122 89171
rect 86178 89115 86246 89171
rect 86302 89115 86326 89171
rect 85726 89047 86326 89115
rect 85726 88991 85750 89047
rect 85806 88991 85874 89047
rect 85930 88991 85998 89047
rect 86054 88991 86122 89047
rect 86178 88991 86246 89047
rect 86302 88991 86326 89047
rect 85726 88923 86326 88991
rect 85726 88867 85750 88923
rect 85806 88867 85874 88923
rect 85930 88867 85998 88923
rect 86054 88867 86122 88923
rect 86178 88867 86246 88923
rect 86302 88867 86326 88923
rect 85726 88799 86326 88867
rect 85726 88743 85750 88799
rect 85806 88743 85874 88799
rect 85930 88743 85998 88799
rect 86054 88743 86122 88799
rect 86178 88743 86246 88799
rect 86302 88743 86326 88799
rect 85726 88675 86326 88743
rect 85726 88619 85750 88675
rect 85806 88619 85874 88675
rect 85930 88619 85998 88675
rect 86054 88619 86122 88675
rect 86178 88619 86246 88675
rect 86302 88619 86326 88675
rect 85726 88551 86326 88619
rect 85726 88495 85750 88551
rect 85806 88495 85874 88551
rect 85930 88495 85998 88551
rect 86054 88495 86122 88551
rect 86178 88495 86246 88551
rect 86302 88495 86326 88551
rect 85726 85889 86326 88495
rect 85726 85833 85750 85889
rect 85806 85833 85874 85889
rect 85930 85833 85998 85889
rect 86054 85833 86122 85889
rect 86178 85833 86246 85889
rect 86302 85833 86326 85889
rect 85726 85765 86326 85833
rect 85726 85709 85750 85765
rect 85806 85709 85874 85765
rect 85930 85709 85998 85765
rect 86054 85709 86122 85765
rect 86178 85709 86246 85765
rect 86302 85709 86326 85765
rect 85726 85641 86326 85709
rect 85726 85585 85750 85641
rect 85806 85585 85874 85641
rect 85930 85585 85998 85641
rect 86054 85585 86122 85641
rect 86178 85585 86246 85641
rect 86302 85585 86326 85641
rect 85726 85517 86326 85585
rect 85726 85461 85750 85517
rect 85806 85461 85874 85517
rect 85930 85461 85998 85517
rect 86054 85461 86122 85517
rect 86178 85461 86246 85517
rect 86302 85461 86326 85517
rect 85726 85393 86326 85461
rect 85726 85337 85750 85393
rect 85806 85337 85874 85393
rect 85930 85337 85998 85393
rect 86054 85337 86122 85393
rect 86178 85337 86246 85393
rect 86302 85337 86326 85393
rect 85726 85269 86326 85337
rect 85726 85213 85750 85269
rect 85806 85213 85874 85269
rect 85930 85213 85998 85269
rect 86054 85213 86122 85269
rect 86178 85213 86246 85269
rect 86302 85213 86326 85269
rect 85726 85145 86326 85213
rect 85726 85089 85750 85145
rect 85806 85089 85874 85145
rect 85930 85089 85998 85145
rect 86054 85089 86122 85145
rect 86178 85089 86246 85145
rect 86302 85089 86326 85145
rect 85726 85021 86326 85089
rect 85726 84965 85750 85021
rect 85806 84965 85874 85021
rect 85930 84965 85998 85021
rect 86054 84965 86122 85021
rect 86178 84965 86246 85021
rect 86302 84965 86326 85021
rect 85726 84897 86326 84965
rect 85726 84841 85750 84897
rect 85806 84841 85874 84897
rect 85930 84841 85998 84897
rect 86054 84841 86122 84897
rect 86178 84841 86246 84897
rect 86302 84841 86326 84897
rect 85726 84773 86326 84841
rect 85726 84717 85750 84773
rect 85806 84717 85874 84773
rect 85930 84717 85998 84773
rect 86054 84717 86122 84773
rect 86178 84717 86246 84773
rect 86302 84717 86326 84773
rect 85726 84649 86326 84717
rect 85726 84593 85750 84649
rect 85806 84593 85874 84649
rect 85930 84593 85998 84649
rect 86054 84593 86122 84649
rect 86178 84593 86246 84649
rect 86302 84593 86326 84649
rect 85726 84525 86326 84593
rect 85726 84469 85750 84525
rect 85806 84469 85874 84525
rect 85930 84469 85998 84525
rect 86054 84469 86122 84525
rect 86178 84469 86246 84525
rect 86302 84469 86326 84525
rect 85726 84401 86326 84469
rect 85726 84345 85750 84401
rect 85806 84345 85874 84401
rect 85930 84345 85998 84401
rect 86054 84345 86122 84401
rect 86178 84345 86246 84401
rect 86302 84345 86326 84401
rect 85726 84277 86326 84345
rect 85726 84221 85750 84277
rect 85806 84221 85874 84277
rect 85930 84221 85998 84277
rect 86054 84221 86122 84277
rect 86178 84221 86246 84277
rect 86302 84221 86326 84277
rect 85726 84153 86326 84221
rect 85726 84097 85750 84153
rect 85806 84097 85874 84153
rect 85930 84097 85998 84153
rect 86054 84097 86122 84153
rect 86178 84097 86246 84153
rect 86302 84097 86326 84153
rect 85726 84029 86326 84097
rect 85726 83973 85750 84029
rect 85806 83973 85874 84029
rect 85930 83973 85998 84029
rect 86054 83973 86122 84029
rect 86178 83973 86246 84029
rect 86302 83973 86326 84029
rect 85726 83905 86326 83973
rect 85726 83849 85750 83905
rect 85806 83849 85874 83905
rect 85930 83849 85998 83905
rect 86054 83849 86122 83905
rect 86178 83849 86246 83905
rect 86302 83849 86326 83905
rect 85726 75000 86326 83849
rect 85726 74944 85750 75000
rect 85806 74944 85874 75000
rect 85930 74944 85998 75000
rect 86054 74944 86122 75000
rect 86178 74944 86246 75000
rect 86302 74944 86326 75000
rect 85726 74876 86326 74944
rect 85726 74820 85750 74876
rect 85806 74820 85874 74876
rect 85930 74820 85998 74876
rect 86054 74820 86122 74876
rect 86178 74820 86246 74876
rect 86302 74820 86326 74876
rect 85726 74752 86326 74820
rect 85726 74696 85750 74752
rect 85806 74696 85874 74752
rect 85930 74696 85998 74752
rect 86054 74696 86122 74752
rect 86178 74696 86246 74752
rect 86302 74696 86326 74752
rect 85726 74628 86326 74696
rect 85726 74572 85750 74628
rect 85806 74572 85874 74628
rect 85930 74572 85998 74628
rect 86054 74572 86122 74628
rect 86178 74572 86246 74628
rect 86302 74572 86326 74628
rect 85726 74504 86326 74572
rect 85726 74448 85750 74504
rect 85806 74448 85874 74504
rect 85930 74448 85998 74504
rect 86054 74448 86122 74504
rect 86178 74448 86246 74504
rect 86302 74448 86326 74504
rect 85726 74380 86326 74448
rect 85726 74324 85750 74380
rect 85806 74324 85874 74380
rect 85930 74324 85998 74380
rect 86054 74324 86122 74380
rect 86178 74324 86246 74380
rect 86302 74324 86326 74380
rect 85726 74256 86326 74324
rect 85726 74200 85750 74256
rect 85806 74200 85874 74256
rect 85930 74200 85998 74256
rect 86054 74200 86122 74256
rect 86178 74200 86246 74256
rect 86302 74200 86326 74256
rect 85726 74132 86326 74200
rect 85726 74076 85750 74132
rect 85806 74076 85874 74132
rect 85930 74076 85998 74132
rect 86054 74076 86122 74132
rect 86178 74076 86246 74132
rect 86302 74076 86326 74132
rect 85726 62064 86326 74076
rect 85726 62008 85812 62064
rect 85868 62008 85936 62064
rect 85992 62008 86060 62064
rect 86116 62008 86184 62064
rect 86240 62008 86326 62064
rect 85726 61940 86326 62008
rect 85726 61884 85812 61940
rect 85868 61884 85936 61940
rect 85992 61884 86060 61940
rect 86116 61884 86184 61940
rect 86240 61884 86326 61940
rect 85726 61816 86326 61884
rect 85726 61760 85812 61816
rect 85868 61760 85936 61816
rect 85992 61760 86060 61816
rect 86116 61760 86184 61816
rect 86240 61760 86326 61816
rect 85726 61692 86326 61760
rect 85726 61636 85812 61692
rect 85868 61636 85936 61692
rect 85992 61636 86060 61692
rect 86116 61636 86184 61692
rect 86240 61636 86326 61692
rect 85726 60264 86326 61636
rect 85726 60208 85812 60264
rect 85868 60208 85936 60264
rect 85992 60208 86060 60264
rect 86116 60208 86184 60264
rect 86240 60208 86326 60264
rect 85726 60140 86326 60208
rect 85726 60084 85812 60140
rect 85868 60084 85936 60140
rect 85992 60084 86060 60140
rect 86116 60084 86184 60140
rect 86240 60084 86326 60140
rect 85726 60016 86326 60084
rect 85726 59960 85812 60016
rect 85868 59960 85936 60016
rect 85992 59960 86060 60016
rect 86116 59960 86184 60016
rect 86240 59960 86326 60016
rect 85726 59892 86326 59960
rect 85726 59836 85812 59892
rect 85868 59836 85936 59892
rect 85992 59836 86060 59892
rect 86116 59836 86184 59892
rect 86240 59836 86326 59892
rect 85726 58464 86326 59836
rect 85726 58408 85812 58464
rect 85868 58408 85936 58464
rect 85992 58408 86060 58464
rect 86116 58408 86184 58464
rect 86240 58408 86326 58464
rect 85726 58340 86326 58408
rect 85726 58284 85812 58340
rect 85868 58284 85936 58340
rect 85992 58284 86060 58340
rect 86116 58284 86184 58340
rect 86240 58284 86326 58340
rect 85726 58216 86326 58284
rect 85726 58160 85812 58216
rect 85868 58160 85936 58216
rect 85992 58160 86060 58216
rect 86116 58160 86184 58216
rect 86240 58160 86326 58216
rect 85726 58092 86326 58160
rect 85726 58036 85812 58092
rect 85868 58036 85936 58092
rect 85992 58036 86060 58092
rect 86116 58036 86184 58092
rect 86240 58036 86326 58092
rect 85726 56664 86326 58036
rect 85726 56608 85812 56664
rect 85868 56608 85936 56664
rect 85992 56608 86060 56664
rect 86116 56608 86184 56664
rect 86240 56608 86326 56664
rect 85726 56540 86326 56608
rect 85726 56484 85812 56540
rect 85868 56484 85936 56540
rect 85992 56484 86060 56540
rect 86116 56484 86184 56540
rect 86240 56484 86326 56540
rect 85726 56416 86326 56484
rect 85726 56360 85812 56416
rect 85868 56360 85936 56416
rect 85992 56360 86060 56416
rect 86116 56360 86184 56416
rect 86240 56360 86326 56416
rect 85726 56292 86326 56360
rect 85726 56236 85812 56292
rect 85868 56236 85936 56292
rect 85992 56236 86060 56292
rect 86116 56236 86184 56292
rect 86240 56236 86326 56292
rect 85726 54864 86326 56236
rect 85726 54808 85812 54864
rect 85868 54808 85936 54864
rect 85992 54808 86060 54864
rect 86116 54808 86184 54864
rect 86240 54808 86326 54864
rect 85726 54740 86326 54808
rect 85726 54684 85812 54740
rect 85868 54684 85936 54740
rect 85992 54684 86060 54740
rect 86116 54684 86184 54740
rect 86240 54684 86326 54740
rect 85726 54616 86326 54684
rect 85726 54560 85812 54616
rect 85868 54560 85936 54616
rect 85992 54560 86060 54616
rect 86116 54560 86184 54616
rect 86240 54560 86326 54616
rect 85726 54492 86326 54560
rect 85726 54436 85812 54492
rect 85868 54436 85936 54492
rect 85992 54436 86060 54492
rect 86116 54436 86184 54492
rect 86240 54436 86326 54492
rect 85726 53064 86326 54436
rect 85726 53008 85812 53064
rect 85868 53008 85936 53064
rect 85992 53008 86060 53064
rect 86116 53008 86184 53064
rect 86240 53008 86326 53064
rect 85726 52940 86326 53008
rect 85726 52884 85812 52940
rect 85868 52884 85936 52940
rect 85992 52884 86060 52940
rect 86116 52884 86184 52940
rect 86240 52884 86326 52940
rect 85726 52816 86326 52884
rect 85726 52760 85812 52816
rect 85868 52760 85936 52816
rect 85992 52760 86060 52816
rect 86116 52760 86184 52816
rect 86240 52760 86326 52816
rect 85726 52692 86326 52760
rect 85726 52636 85812 52692
rect 85868 52636 85936 52692
rect 85992 52636 86060 52692
rect 86116 52636 86184 52692
rect 86240 52636 86326 52692
rect 85726 51264 86326 52636
rect 85726 51208 85812 51264
rect 85868 51208 85936 51264
rect 85992 51208 86060 51264
rect 86116 51208 86184 51264
rect 86240 51208 86326 51264
rect 85726 51140 86326 51208
rect 85726 51084 85812 51140
rect 85868 51084 85936 51140
rect 85992 51084 86060 51140
rect 86116 51084 86184 51140
rect 86240 51084 86326 51140
rect 85726 51016 86326 51084
rect 85726 50960 85812 51016
rect 85868 50960 85936 51016
rect 85992 50960 86060 51016
rect 86116 50960 86184 51016
rect 86240 50960 86326 51016
rect 85726 50892 86326 50960
rect 85726 50836 85812 50892
rect 85868 50836 85936 50892
rect 85992 50836 86060 50892
rect 86116 50836 86184 50892
rect 86240 50836 86326 50892
rect 85726 49464 86326 50836
rect 85726 49408 85812 49464
rect 85868 49408 85936 49464
rect 85992 49408 86060 49464
rect 86116 49408 86184 49464
rect 86240 49408 86326 49464
rect 85726 49340 86326 49408
rect 85726 49284 85812 49340
rect 85868 49284 85936 49340
rect 85992 49284 86060 49340
rect 86116 49284 86184 49340
rect 86240 49284 86326 49340
rect 85726 49216 86326 49284
rect 85726 49160 85812 49216
rect 85868 49160 85936 49216
rect 85992 49160 86060 49216
rect 86116 49160 86184 49216
rect 86240 49160 86326 49216
rect 85726 49092 86326 49160
rect 85726 49036 85812 49092
rect 85868 49036 85936 49092
rect 85992 49036 86060 49092
rect 86116 49036 86184 49092
rect 86240 49036 86326 49092
rect 85726 47664 86326 49036
rect 85726 47608 85812 47664
rect 85868 47608 85936 47664
rect 85992 47608 86060 47664
rect 86116 47608 86184 47664
rect 86240 47608 86326 47664
rect 85726 47540 86326 47608
rect 85726 47484 85812 47540
rect 85868 47484 85936 47540
rect 85992 47484 86060 47540
rect 86116 47484 86184 47540
rect 86240 47484 86326 47540
rect 85726 47416 86326 47484
rect 85726 47360 85812 47416
rect 85868 47360 85936 47416
rect 85992 47360 86060 47416
rect 86116 47360 86184 47416
rect 86240 47360 86326 47416
rect 85726 47292 86326 47360
rect 85726 47236 85812 47292
rect 85868 47236 85936 47292
rect 85992 47236 86060 47292
rect 86116 47236 86184 47292
rect 86240 47236 86326 47292
rect 85726 45864 86326 47236
rect 85726 45808 85812 45864
rect 85868 45808 85936 45864
rect 85992 45808 86060 45864
rect 86116 45808 86184 45864
rect 86240 45808 86326 45864
rect 85726 45740 86326 45808
rect 85726 45684 85812 45740
rect 85868 45684 85936 45740
rect 85992 45684 86060 45740
rect 86116 45684 86184 45740
rect 86240 45684 86326 45740
rect 85726 45616 86326 45684
rect 85726 45560 85812 45616
rect 85868 45560 85936 45616
rect 85992 45560 86060 45616
rect 86116 45560 86184 45616
rect 86240 45560 86326 45616
rect 85726 45492 86326 45560
rect 85726 45436 85812 45492
rect 85868 45436 85936 45492
rect 85992 45436 86060 45492
rect 86116 45436 86184 45492
rect 86240 45436 86326 45492
rect 85726 44064 86326 45436
rect 85726 44008 85812 44064
rect 85868 44008 85936 44064
rect 85992 44008 86060 44064
rect 86116 44008 86184 44064
rect 86240 44008 86326 44064
rect 85726 43940 86326 44008
rect 85726 43884 85812 43940
rect 85868 43884 85936 43940
rect 85992 43884 86060 43940
rect 86116 43884 86184 43940
rect 86240 43884 86326 43940
rect 85726 43816 86326 43884
rect 85726 43760 85812 43816
rect 85868 43760 85936 43816
rect 85992 43760 86060 43816
rect 86116 43760 86184 43816
rect 86240 43760 86326 43816
rect 85726 43692 86326 43760
rect 85726 43636 85812 43692
rect 85868 43636 85936 43692
rect 85992 43636 86060 43692
rect 86116 43636 86184 43692
rect 86240 43636 86326 43692
rect 85726 42264 86326 43636
rect 85726 42208 85812 42264
rect 85868 42208 85936 42264
rect 85992 42208 86060 42264
rect 86116 42208 86184 42264
rect 86240 42208 86326 42264
rect 85726 42140 86326 42208
rect 85726 42084 85812 42140
rect 85868 42084 85936 42140
rect 85992 42084 86060 42140
rect 86116 42084 86184 42140
rect 86240 42084 86326 42140
rect 85726 42016 86326 42084
rect 85726 41960 85812 42016
rect 85868 41960 85936 42016
rect 85992 41960 86060 42016
rect 86116 41960 86184 42016
rect 86240 41960 86326 42016
rect 85726 41892 86326 41960
rect 85726 41836 85812 41892
rect 85868 41836 85936 41892
rect 85992 41836 86060 41892
rect 86116 41836 86184 41892
rect 86240 41836 86326 41892
rect 85726 40464 86326 41836
rect 85726 40408 85812 40464
rect 85868 40408 85936 40464
rect 85992 40408 86060 40464
rect 86116 40408 86184 40464
rect 86240 40408 86326 40464
rect 85726 40340 86326 40408
rect 85726 40284 85812 40340
rect 85868 40284 85936 40340
rect 85992 40284 86060 40340
rect 86116 40284 86184 40340
rect 86240 40284 86326 40340
rect 85726 40216 86326 40284
rect 85726 40160 85812 40216
rect 85868 40160 85936 40216
rect 85992 40160 86060 40216
rect 86116 40160 86184 40216
rect 86240 40160 86326 40216
rect 85726 40092 86326 40160
rect 85726 40036 85812 40092
rect 85868 40036 85936 40092
rect 85992 40036 86060 40092
rect 86116 40036 86184 40092
rect 86240 40036 86326 40092
rect 85726 38664 86326 40036
rect 85726 38608 85812 38664
rect 85868 38608 85936 38664
rect 85992 38608 86060 38664
rect 86116 38608 86184 38664
rect 86240 38608 86326 38664
rect 85726 38540 86326 38608
rect 85726 38484 85812 38540
rect 85868 38484 85936 38540
rect 85992 38484 86060 38540
rect 86116 38484 86184 38540
rect 86240 38484 86326 38540
rect 85726 38416 86326 38484
rect 85726 38360 85812 38416
rect 85868 38360 85936 38416
rect 85992 38360 86060 38416
rect 86116 38360 86184 38416
rect 86240 38360 86326 38416
rect 85726 38292 86326 38360
rect 85726 38236 85812 38292
rect 85868 38236 85936 38292
rect 85992 38236 86060 38292
rect 86116 38236 86184 38292
rect 86240 38236 86326 38292
rect 85726 36864 86326 38236
rect 85726 36808 85812 36864
rect 85868 36808 85936 36864
rect 85992 36808 86060 36864
rect 86116 36808 86184 36864
rect 86240 36808 86326 36864
rect 85726 36740 86326 36808
rect 85726 36684 85812 36740
rect 85868 36684 85936 36740
rect 85992 36684 86060 36740
rect 86116 36684 86184 36740
rect 86240 36684 86326 36740
rect 85726 36616 86326 36684
rect 85726 36560 85812 36616
rect 85868 36560 85936 36616
rect 85992 36560 86060 36616
rect 86116 36560 86184 36616
rect 86240 36560 86326 36616
rect 85726 36492 86326 36560
rect 85726 36436 85812 36492
rect 85868 36436 85936 36492
rect 85992 36436 86060 36492
rect 86116 36436 86184 36492
rect 86240 36436 86326 36492
rect 85726 35064 86326 36436
rect 85726 35008 85812 35064
rect 85868 35008 85936 35064
rect 85992 35008 86060 35064
rect 86116 35008 86184 35064
rect 86240 35008 86326 35064
rect 85726 34940 86326 35008
rect 85726 34884 85812 34940
rect 85868 34884 85936 34940
rect 85992 34884 86060 34940
rect 86116 34884 86184 34940
rect 86240 34884 86326 34940
rect 85726 34816 86326 34884
rect 85726 34760 85812 34816
rect 85868 34760 85936 34816
rect 85992 34760 86060 34816
rect 86116 34760 86184 34816
rect 86240 34760 86326 34816
rect 85726 34692 86326 34760
rect 85726 34636 85812 34692
rect 85868 34636 85936 34692
rect 85992 34636 86060 34692
rect 86116 34636 86184 34692
rect 86240 34636 86326 34692
rect 85726 33264 86326 34636
rect 85726 33208 85812 33264
rect 85868 33208 85936 33264
rect 85992 33208 86060 33264
rect 86116 33208 86184 33264
rect 86240 33208 86326 33264
rect 85726 33140 86326 33208
rect 85726 33084 85812 33140
rect 85868 33084 85936 33140
rect 85992 33084 86060 33140
rect 86116 33084 86184 33140
rect 86240 33084 86326 33140
rect 85726 33016 86326 33084
rect 85726 32960 85812 33016
rect 85868 32960 85936 33016
rect 85992 32960 86060 33016
rect 86116 32960 86184 33016
rect 86240 32960 86326 33016
rect 85726 32892 86326 32960
rect 85726 32836 85812 32892
rect 85868 32836 85936 32892
rect 85992 32836 86060 32892
rect 86116 32836 86184 32892
rect 86240 32836 86326 32892
rect 85726 31464 86326 32836
rect 85726 31408 85812 31464
rect 85868 31408 85936 31464
rect 85992 31408 86060 31464
rect 86116 31408 86184 31464
rect 86240 31408 86326 31464
rect 85726 31340 86326 31408
rect 85726 31284 85812 31340
rect 85868 31284 85936 31340
rect 85992 31284 86060 31340
rect 86116 31284 86184 31340
rect 86240 31284 86326 31340
rect 85726 31216 86326 31284
rect 85726 31160 85812 31216
rect 85868 31160 85936 31216
rect 85992 31160 86060 31216
rect 86116 31160 86184 31216
rect 86240 31160 86326 31216
rect 85726 31092 86326 31160
rect 85726 31036 85812 31092
rect 85868 31036 85936 31092
rect 85992 31036 86060 31092
rect 86116 31036 86184 31092
rect 86240 31036 86326 31092
rect 85726 29664 86326 31036
rect 85726 29608 85812 29664
rect 85868 29608 85936 29664
rect 85992 29608 86060 29664
rect 86116 29608 86184 29664
rect 86240 29608 86326 29664
rect 85726 29540 86326 29608
rect 85726 29484 85812 29540
rect 85868 29484 85936 29540
rect 85992 29484 86060 29540
rect 86116 29484 86184 29540
rect 86240 29484 86326 29540
rect 85726 29416 86326 29484
rect 85726 29360 85812 29416
rect 85868 29360 85936 29416
rect 85992 29360 86060 29416
rect 86116 29360 86184 29416
rect 86240 29360 86326 29416
rect 85726 29292 86326 29360
rect 85726 29236 85812 29292
rect 85868 29236 85936 29292
rect 85992 29236 86060 29292
rect 86116 29236 86184 29292
rect 86240 29236 86326 29292
rect 85726 27864 86326 29236
rect 85726 27808 85812 27864
rect 85868 27808 85936 27864
rect 85992 27808 86060 27864
rect 86116 27808 86184 27864
rect 86240 27808 86326 27864
rect 85726 27740 86326 27808
rect 85726 27684 85812 27740
rect 85868 27684 85936 27740
rect 85992 27684 86060 27740
rect 86116 27684 86184 27740
rect 86240 27684 86326 27740
rect 85726 27616 86326 27684
rect 85726 27560 85812 27616
rect 85868 27560 85936 27616
rect 85992 27560 86060 27616
rect 86116 27560 86184 27616
rect 86240 27560 86326 27616
rect 85726 27492 86326 27560
rect 85726 27436 85812 27492
rect 85868 27436 85936 27492
rect 85992 27436 86060 27492
rect 86116 27436 86184 27492
rect 86240 27436 86326 27492
rect 85726 26064 86326 27436
rect 85726 26008 85812 26064
rect 85868 26008 85936 26064
rect 85992 26008 86060 26064
rect 86116 26008 86184 26064
rect 86240 26008 86326 26064
rect 85726 25940 86326 26008
rect 85726 25884 85812 25940
rect 85868 25884 85936 25940
rect 85992 25884 86060 25940
rect 86116 25884 86184 25940
rect 86240 25884 86326 25940
rect 85726 25816 86326 25884
rect 85726 25760 85812 25816
rect 85868 25760 85936 25816
rect 85992 25760 86060 25816
rect 86116 25760 86184 25816
rect 86240 25760 86326 25816
rect 85726 25692 86326 25760
rect 85726 25636 85812 25692
rect 85868 25636 85936 25692
rect 85992 25636 86060 25692
rect 86116 25636 86184 25692
rect 86240 25636 86326 25692
rect 85726 24264 86326 25636
rect 85726 24208 85812 24264
rect 85868 24208 85936 24264
rect 85992 24208 86060 24264
rect 86116 24208 86184 24264
rect 86240 24208 86326 24264
rect 85726 24140 86326 24208
rect 85726 24084 85812 24140
rect 85868 24084 85936 24140
rect 85992 24084 86060 24140
rect 86116 24084 86184 24140
rect 86240 24084 86326 24140
rect 85726 24016 86326 24084
rect 85726 23960 85812 24016
rect 85868 23960 85936 24016
rect 85992 23960 86060 24016
rect 86116 23960 86184 24016
rect 86240 23960 86326 24016
rect 85726 23892 86326 23960
rect 85726 23836 85812 23892
rect 85868 23836 85936 23892
rect 85992 23836 86060 23892
rect 86116 23836 86184 23892
rect 86240 23836 86326 23892
rect 85726 22464 86326 23836
rect 85726 22408 85812 22464
rect 85868 22408 85936 22464
rect 85992 22408 86060 22464
rect 86116 22408 86184 22464
rect 86240 22408 86326 22464
rect 85726 22340 86326 22408
rect 85726 22284 85812 22340
rect 85868 22284 85936 22340
rect 85992 22284 86060 22340
rect 86116 22284 86184 22340
rect 86240 22284 86326 22340
rect 85726 22216 86326 22284
rect 85726 22160 85812 22216
rect 85868 22160 85936 22216
rect 85992 22160 86060 22216
rect 86116 22160 86184 22216
rect 86240 22160 86326 22216
rect 85726 22092 86326 22160
rect 85726 22036 85812 22092
rect 85868 22036 85936 22092
rect 85992 22036 86060 22092
rect 86116 22036 86184 22092
rect 86240 22036 86326 22092
rect 85726 20664 86326 22036
rect 85726 20608 85812 20664
rect 85868 20608 85936 20664
rect 85992 20608 86060 20664
rect 86116 20608 86184 20664
rect 86240 20608 86326 20664
rect 85726 20540 86326 20608
rect 85726 20484 85812 20540
rect 85868 20484 85936 20540
rect 85992 20484 86060 20540
rect 86116 20484 86184 20540
rect 86240 20484 86326 20540
rect 85726 20416 86326 20484
rect 85726 20360 85812 20416
rect 85868 20360 85936 20416
rect 85992 20360 86060 20416
rect 86116 20360 86184 20416
rect 86240 20360 86326 20416
rect 85726 20292 86326 20360
rect 85726 20236 85812 20292
rect 85868 20236 85936 20292
rect 85992 20236 86060 20292
rect 86116 20236 86184 20292
rect 86240 20236 86326 20292
rect 85726 18864 86326 20236
rect 85726 18808 85812 18864
rect 85868 18808 85936 18864
rect 85992 18808 86060 18864
rect 86116 18808 86184 18864
rect 86240 18808 86326 18864
rect 85726 18740 86326 18808
rect 85726 18684 85812 18740
rect 85868 18684 85936 18740
rect 85992 18684 86060 18740
rect 86116 18684 86184 18740
rect 86240 18684 86326 18740
rect 85726 18616 86326 18684
rect 85726 18560 85812 18616
rect 85868 18560 85936 18616
rect 85992 18560 86060 18616
rect 86116 18560 86184 18616
rect 86240 18560 86326 18616
rect 85726 18492 86326 18560
rect 85726 18436 85812 18492
rect 85868 18436 85936 18492
rect 85992 18436 86060 18492
rect 86116 18436 86184 18492
rect 86240 18436 86326 18492
rect 85726 17064 86326 18436
rect 85726 17008 85812 17064
rect 85868 17008 85936 17064
rect 85992 17008 86060 17064
rect 86116 17008 86184 17064
rect 86240 17008 86326 17064
rect 85726 16940 86326 17008
rect 85726 16884 85812 16940
rect 85868 16884 85936 16940
rect 85992 16884 86060 16940
rect 86116 16884 86184 16940
rect 86240 16884 86326 16940
rect 85726 16816 86326 16884
rect 85726 16760 85812 16816
rect 85868 16760 85936 16816
rect 85992 16760 86060 16816
rect 86116 16760 86184 16816
rect 86240 16760 86326 16816
rect 85726 16692 86326 16760
rect 85726 16636 85812 16692
rect 85868 16636 85936 16692
rect 85992 16636 86060 16692
rect 86116 16636 86184 16692
rect 86240 16636 86326 16692
rect 85726 15264 86326 16636
rect 85726 15208 85812 15264
rect 85868 15208 85936 15264
rect 85992 15208 86060 15264
rect 86116 15208 86184 15264
rect 86240 15208 86326 15264
rect 85726 15140 86326 15208
rect 85726 15084 85812 15140
rect 85868 15084 85936 15140
rect 85992 15084 86060 15140
rect 86116 15084 86184 15140
rect 86240 15084 86326 15140
rect 85726 15016 86326 15084
rect 85726 14960 85812 15016
rect 85868 14960 85936 15016
rect 85992 14960 86060 15016
rect 86116 14960 86184 15016
rect 86240 14960 86326 15016
rect 85726 14892 86326 14960
rect 85726 14836 85812 14892
rect 85868 14836 85936 14892
rect 85992 14836 86060 14892
rect 86116 14836 86184 14892
rect 86240 14836 86326 14892
rect 85726 13464 86326 14836
rect 85726 13408 85812 13464
rect 85868 13408 85936 13464
rect 85992 13408 86060 13464
rect 86116 13408 86184 13464
rect 86240 13408 86326 13464
rect 85726 13340 86326 13408
rect 85726 13284 85812 13340
rect 85868 13284 85936 13340
rect 85992 13284 86060 13340
rect 86116 13284 86184 13340
rect 86240 13284 86326 13340
rect 85726 13216 86326 13284
rect 85726 13160 85812 13216
rect 85868 13160 85936 13216
rect 85992 13160 86060 13216
rect 86116 13160 86184 13216
rect 86240 13160 86326 13216
rect 85726 13092 86326 13160
rect 85726 13036 85812 13092
rect 85868 13036 85936 13092
rect 85992 13036 86060 13092
rect 86116 13036 86184 13092
rect 86240 13036 86326 13092
rect 85726 11664 86326 13036
rect 85726 11608 85812 11664
rect 85868 11608 85936 11664
rect 85992 11608 86060 11664
rect 86116 11608 86184 11664
rect 86240 11608 86326 11664
rect 85726 11540 86326 11608
rect 85726 11484 85812 11540
rect 85868 11484 85936 11540
rect 85992 11484 86060 11540
rect 86116 11484 86184 11540
rect 86240 11484 86326 11540
rect 85726 11416 86326 11484
rect 85726 11360 85812 11416
rect 85868 11360 85936 11416
rect 85992 11360 86060 11416
rect 86116 11360 86184 11416
rect 86240 11360 86326 11416
rect 85726 11292 86326 11360
rect 85726 11236 85812 11292
rect 85868 11236 85936 11292
rect 85992 11236 86060 11292
rect 86116 11236 86184 11292
rect 86240 11236 86326 11292
rect 85726 9864 86326 11236
rect 85726 9808 85812 9864
rect 85868 9808 85936 9864
rect 85992 9808 86060 9864
rect 86116 9808 86184 9864
rect 86240 9808 86326 9864
rect 85726 9740 86326 9808
rect 85726 9684 85812 9740
rect 85868 9684 85936 9740
rect 85992 9684 86060 9740
rect 86116 9684 86184 9740
rect 86240 9684 86326 9740
rect 85726 9616 86326 9684
rect 85726 9560 85812 9616
rect 85868 9560 85936 9616
rect 85992 9560 86060 9616
rect 86116 9560 86184 9616
rect 86240 9560 86326 9616
rect 85726 9492 86326 9560
rect 85726 9436 85812 9492
rect 85868 9436 85936 9492
rect 85992 9436 86060 9492
rect 86116 9436 86184 9492
rect 86240 9436 86326 9492
rect 85726 8064 86326 9436
rect 85726 8008 85812 8064
rect 85868 8008 85936 8064
rect 85992 8008 86060 8064
rect 86116 8008 86184 8064
rect 86240 8008 86326 8064
rect 85726 7940 86326 8008
rect 85726 7884 85812 7940
rect 85868 7884 85936 7940
rect 85992 7884 86060 7940
rect 86116 7884 86184 7940
rect 86240 7884 86326 7940
rect 85726 7816 86326 7884
rect 85726 7760 85812 7816
rect 85868 7760 85936 7816
rect 85992 7760 86060 7816
rect 86116 7760 86184 7816
rect 86240 7760 86326 7816
rect 85726 7692 86326 7760
rect 85726 7636 85812 7692
rect 85868 7636 85936 7692
rect 85992 7636 86060 7692
rect 86116 7636 86184 7692
rect 86240 7636 86326 7692
rect 85726 6264 86326 7636
rect 85726 6208 85812 6264
rect 85868 6208 85936 6264
rect 85992 6208 86060 6264
rect 86116 6208 86184 6264
rect 86240 6208 86326 6264
rect 85726 6140 86326 6208
rect 85726 6084 85812 6140
rect 85868 6084 85936 6140
rect 85992 6084 86060 6140
rect 86116 6084 86184 6140
rect 86240 6084 86326 6140
rect 85726 6016 86326 6084
rect 85726 5960 85812 6016
rect 85868 5960 85936 6016
rect 85992 5960 86060 6016
rect 86116 5960 86184 6016
rect 86240 5960 86326 6016
rect 85726 5892 86326 5960
rect 85726 5836 85812 5892
rect 85868 5836 85936 5892
rect 85992 5836 86060 5892
rect 86116 5836 86184 5892
rect 86240 5836 86326 5892
rect 85726 4464 86326 5836
rect 85726 4408 85812 4464
rect 85868 4408 85936 4464
rect 85992 4408 86060 4464
rect 86116 4408 86184 4464
rect 86240 4408 86326 4464
rect 85726 4340 86326 4408
rect 85726 4284 85812 4340
rect 85868 4284 85936 4340
rect 85992 4284 86060 4340
rect 86116 4284 86184 4340
rect 86240 4284 86326 4340
rect 85726 4216 86326 4284
rect 85726 4160 85812 4216
rect 85868 4160 85936 4216
rect 85992 4160 86060 4216
rect 86116 4160 86184 4216
rect 86240 4160 86326 4216
rect 85726 4092 86326 4160
rect 85726 4036 85812 4092
rect 85868 4036 85936 4092
rect 85992 4036 86060 4092
rect 86116 4036 86184 4092
rect 86240 4036 86326 4092
rect 85726 3136 86326 4036
rect 86526 95425 87126 95648
rect 86526 95369 86550 95425
rect 86606 95369 86674 95425
rect 86730 95369 86798 95425
rect 86854 95369 86922 95425
rect 86978 95369 87046 95425
rect 87102 95369 87126 95425
rect 86526 95301 87126 95369
rect 86526 95245 86550 95301
rect 86606 95245 86674 95301
rect 86730 95245 86798 95301
rect 86854 95245 86922 95301
rect 86978 95245 87046 95301
rect 87102 95245 87126 95301
rect 86526 95177 87126 95245
rect 86526 95121 86550 95177
rect 86606 95121 86674 95177
rect 86730 95121 86798 95177
rect 86854 95121 86922 95177
rect 86978 95121 87046 95177
rect 87102 95121 87126 95177
rect 86526 95053 87126 95121
rect 86526 94997 86550 95053
rect 86606 94997 86674 95053
rect 86730 94997 86798 95053
rect 86854 94997 86922 95053
rect 86978 94997 87046 95053
rect 87102 94997 87126 95053
rect 86526 94929 87126 94997
rect 86526 94873 86550 94929
rect 86606 94873 86674 94929
rect 86730 94873 86798 94929
rect 86854 94873 86922 94929
rect 86978 94873 87046 94929
rect 87102 94873 87126 94929
rect 86526 94805 87126 94873
rect 86526 94749 86550 94805
rect 86606 94749 86674 94805
rect 86730 94749 86798 94805
rect 86854 94749 86922 94805
rect 86978 94749 87046 94805
rect 87102 94749 87126 94805
rect 86526 94681 87126 94749
rect 86526 94625 86550 94681
rect 86606 94625 86674 94681
rect 86730 94625 86798 94681
rect 86854 94625 86922 94681
rect 86978 94625 87046 94681
rect 87102 94625 87126 94681
rect 86526 94557 87126 94625
rect 86526 94501 86550 94557
rect 86606 94501 86674 94557
rect 86730 94501 86798 94557
rect 86854 94501 86922 94557
rect 86978 94501 87046 94557
rect 87102 94501 87126 94557
rect 86526 94433 87126 94501
rect 86526 94377 86550 94433
rect 86606 94377 86674 94433
rect 86730 94377 86798 94433
rect 86854 94377 86922 94433
rect 86978 94377 87046 94433
rect 87102 94377 87126 94433
rect 86526 94309 87126 94377
rect 86526 94253 86550 94309
rect 86606 94253 86674 94309
rect 86730 94253 86798 94309
rect 86854 94253 86922 94309
rect 86978 94253 87046 94309
rect 87102 94253 87126 94309
rect 86526 92191 87126 94253
rect 86526 92135 86550 92191
rect 86606 92135 86674 92191
rect 86730 92135 86798 92191
rect 86854 92135 86922 92191
rect 86978 92135 87046 92191
rect 87102 92135 87126 92191
rect 86526 92067 87126 92135
rect 86526 92011 86550 92067
rect 86606 92011 86674 92067
rect 86730 92011 86798 92067
rect 86854 92011 86922 92067
rect 86978 92011 87046 92067
rect 87102 92011 87126 92067
rect 86526 91943 87126 92011
rect 86526 91887 86550 91943
rect 86606 91887 86674 91943
rect 86730 91887 86798 91943
rect 86854 91887 86922 91943
rect 86978 91887 87046 91943
rect 87102 91887 87126 91943
rect 86526 91819 87126 91887
rect 86526 91763 86550 91819
rect 86606 91763 86674 91819
rect 86730 91763 86798 91819
rect 86854 91763 86922 91819
rect 86978 91763 87046 91819
rect 87102 91763 87126 91819
rect 86526 91695 87126 91763
rect 86526 91639 86550 91695
rect 86606 91639 86674 91695
rect 86730 91639 86798 91695
rect 86854 91639 86922 91695
rect 86978 91639 87046 91695
rect 87102 91639 87126 91695
rect 86526 91571 87126 91639
rect 86526 91515 86550 91571
rect 86606 91515 86674 91571
rect 86730 91515 86798 91571
rect 86854 91515 86922 91571
rect 86978 91515 87046 91571
rect 87102 91515 87126 91571
rect 86526 91447 87126 91515
rect 86526 91391 86550 91447
rect 86606 91391 86674 91447
rect 86730 91391 86798 91447
rect 86854 91391 86922 91447
rect 86978 91391 87046 91447
rect 87102 91391 87126 91447
rect 86526 91323 87126 91391
rect 86526 91267 86550 91323
rect 86606 91267 86674 91323
rect 86730 91267 86798 91323
rect 86854 91267 86922 91323
rect 86978 91267 87046 91323
rect 87102 91267 87126 91323
rect 86526 91199 87126 91267
rect 86526 91143 86550 91199
rect 86606 91143 86674 91199
rect 86730 91143 86798 91199
rect 86854 91143 86922 91199
rect 86978 91143 87046 91199
rect 87102 91143 87126 91199
rect 86526 91075 87126 91143
rect 86526 91019 86550 91075
rect 86606 91019 86674 91075
rect 86730 91019 86798 91075
rect 86854 91019 86922 91075
rect 86978 91019 87046 91075
rect 87102 91019 87126 91075
rect 86526 90951 87126 91019
rect 86526 90895 86550 90951
rect 86606 90895 86674 90951
rect 86730 90895 86798 90951
rect 86854 90895 86922 90951
rect 86978 90895 87046 90951
rect 87102 90895 87126 90951
rect 86526 90827 87126 90895
rect 86526 90771 86550 90827
rect 86606 90771 86674 90827
rect 86730 90771 86798 90827
rect 86854 90771 86922 90827
rect 86978 90771 87046 90827
rect 87102 90771 87126 90827
rect 86526 90703 87126 90771
rect 86526 90647 86550 90703
rect 86606 90647 86674 90703
rect 86730 90647 86798 90703
rect 86854 90647 86922 90703
rect 86978 90647 87046 90703
rect 87102 90647 87126 90703
rect 86526 90579 87126 90647
rect 86526 90523 86550 90579
rect 86606 90523 86674 90579
rect 86730 90523 86798 90579
rect 86854 90523 86922 90579
rect 86978 90523 87046 90579
rect 87102 90523 87126 90579
rect 86526 90455 87126 90523
rect 86526 90399 86550 90455
rect 86606 90399 86674 90455
rect 86730 90399 86798 90455
rect 86854 90399 86922 90455
rect 86978 90399 87046 90455
rect 87102 90399 87126 90455
rect 86526 83587 87126 90399
rect 86526 83531 86550 83587
rect 86606 83531 86674 83587
rect 86730 83531 86798 83587
rect 86854 83531 86922 83587
rect 86978 83531 87046 83587
rect 87102 83531 87126 83587
rect 86526 83463 87126 83531
rect 86526 83407 86550 83463
rect 86606 83407 86674 83463
rect 86730 83407 86798 83463
rect 86854 83407 86922 83463
rect 86978 83407 87046 83463
rect 87102 83407 87126 83463
rect 86526 83339 87126 83407
rect 86526 83283 86550 83339
rect 86606 83283 86674 83339
rect 86730 83283 86798 83339
rect 86854 83283 86922 83339
rect 86978 83283 87046 83339
rect 87102 83283 87126 83339
rect 86526 83215 87126 83283
rect 86526 83159 86550 83215
rect 86606 83159 86674 83215
rect 86730 83159 86798 83215
rect 86854 83159 86922 83215
rect 86978 83159 87046 83215
rect 87102 83159 87126 83215
rect 86526 83091 87126 83159
rect 86526 83035 86550 83091
rect 86606 83035 86674 83091
rect 86730 83035 86798 83091
rect 86854 83035 86922 83091
rect 86978 83035 87046 83091
rect 87102 83035 87126 83091
rect 86526 82967 87126 83035
rect 86526 82911 86550 82967
rect 86606 82911 86674 82967
rect 86730 82911 86798 82967
rect 86854 82911 86922 82967
rect 86978 82911 87046 82967
rect 87102 82911 87126 82967
rect 86526 82843 87126 82911
rect 86526 82787 86550 82843
rect 86606 82787 86674 82843
rect 86730 82787 86798 82843
rect 86854 82787 86922 82843
rect 86978 82787 87046 82843
rect 87102 82787 87126 82843
rect 86526 82719 87126 82787
rect 86526 82663 86550 82719
rect 86606 82663 86674 82719
rect 86730 82663 86798 82719
rect 86854 82663 86922 82719
rect 86978 82663 87046 82719
rect 87102 82663 87126 82719
rect 86526 82595 87126 82663
rect 86526 82539 86550 82595
rect 86606 82539 86674 82595
rect 86730 82539 86798 82595
rect 86854 82539 86922 82595
rect 86978 82539 87046 82595
rect 87102 82539 87126 82595
rect 86526 82471 87126 82539
rect 86526 82415 86550 82471
rect 86606 82415 86674 82471
rect 86730 82415 86798 82471
rect 86854 82415 86922 82471
rect 86978 82415 87046 82471
rect 87102 82415 87126 82471
rect 86526 82347 87126 82415
rect 86526 82291 86550 82347
rect 86606 82291 86674 82347
rect 86730 82291 86798 82347
rect 86854 82291 86922 82347
rect 86978 82291 87046 82347
rect 87102 82291 87126 82347
rect 86526 82223 87126 82291
rect 86526 82167 86550 82223
rect 86606 82167 86674 82223
rect 86730 82167 86798 82223
rect 86854 82167 86922 82223
rect 86978 82167 87046 82223
rect 87102 82167 87126 82223
rect 86526 82099 87126 82167
rect 86526 82043 86550 82099
rect 86606 82043 86674 82099
rect 86730 82043 86798 82099
rect 86854 82043 86922 82099
rect 86978 82043 87046 82099
rect 87102 82043 87126 82099
rect 86526 81975 87126 82043
rect 86526 81919 86550 81975
rect 86606 81919 86674 81975
rect 86730 81919 86798 81975
rect 86854 81919 86922 81975
rect 86978 81919 87046 81975
rect 87102 81919 87126 81975
rect 86526 81851 87126 81919
rect 86526 81795 86550 81851
rect 86606 81795 86674 81851
rect 86730 81795 86798 81851
rect 86854 81795 86922 81851
rect 86978 81795 87046 81851
rect 87102 81795 87126 81851
rect 86526 81727 87126 81795
rect 86526 81671 86550 81727
rect 86606 81671 86674 81727
rect 86730 81671 86798 81727
rect 86854 81671 86922 81727
rect 86978 81671 87046 81727
rect 87102 81671 87126 81727
rect 86526 81603 87126 81671
rect 86526 81547 86550 81603
rect 86606 81547 86674 81603
rect 86730 81547 86798 81603
rect 86854 81547 86922 81603
rect 86978 81547 87046 81603
rect 87102 81547 87126 81603
rect 86526 81479 87126 81547
rect 86526 81423 86550 81479
rect 86606 81423 86674 81479
rect 86730 81423 86798 81479
rect 86854 81423 86922 81479
rect 86978 81423 87046 81479
rect 87102 81423 87126 81479
rect 86526 81355 87126 81423
rect 86526 81299 86550 81355
rect 86606 81299 86674 81355
rect 86730 81299 86798 81355
rect 86854 81299 86922 81355
rect 86978 81299 87046 81355
rect 87102 81299 87126 81355
rect 86526 81231 87126 81299
rect 86526 81175 86550 81231
rect 86606 81175 86674 81231
rect 86730 81175 86798 81231
rect 86854 81175 86922 81231
rect 86978 81175 87046 81231
rect 87102 81175 87126 81231
rect 86526 81107 87126 81175
rect 86526 81051 86550 81107
rect 86606 81051 86674 81107
rect 86730 81051 86798 81107
rect 86854 81051 86922 81107
rect 86978 81051 87046 81107
rect 87102 81051 87126 81107
rect 86526 80983 87126 81051
rect 86526 80927 86550 80983
rect 86606 80927 86674 80983
rect 86730 80927 86798 80983
rect 86854 80927 86922 80983
rect 86978 80927 87046 80983
rect 87102 80927 87126 80983
rect 86526 80859 87126 80927
rect 86526 80803 86550 80859
rect 86606 80803 86674 80859
rect 86730 80803 86798 80859
rect 86854 80803 86922 80859
rect 86978 80803 87046 80859
rect 87102 80803 87126 80859
rect 86526 80735 87126 80803
rect 86526 80679 86550 80735
rect 86606 80679 86674 80735
rect 86730 80679 86798 80735
rect 86854 80679 86922 80735
rect 86978 80679 87046 80735
rect 87102 80679 87126 80735
rect 86526 80611 87126 80679
rect 86526 80555 86550 80611
rect 86606 80555 86674 80611
rect 86730 80555 86798 80611
rect 86854 80555 86922 80611
rect 86978 80555 87046 80611
rect 87102 80555 87126 80611
rect 86526 80487 87126 80555
rect 86526 80431 86550 80487
rect 86606 80431 86674 80487
rect 86730 80431 86798 80487
rect 86854 80431 86922 80487
rect 86978 80431 87046 80487
rect 87102 80431 87126 80487
rect 86526 80363 87126 80431
rect 86526 80307 86550 80363
rect 86606 80307 86674 80363
rect 86730 80307 86798 80363
rect 86854 80307 86922 80363
rect 86978 80307 87046 80363
rect 87102 80307 87126 80363
rect 86526 76656 87126 80307
rect 86526 76600 86550 76656
rect 86606 76600 86674 76656
rect 86730 76600 86798 76656
rect 86854 76600 86922 76656
rect 86978 76600 87046 76656
rect 87102 76600 87126 76656
rect 86526 76532 87126 76600
rect 86526 76476 86550 76532
rect 86606 76476 86674 76532
rect 86730 76476 86798 76532
rect 86854 76476 86922 76532
rect 86978 76476 87046 76532
rect 87102 76476 87126 76532
rect 86526 76408 87126 76476
rect 86526 76352 86550 76408
rect 86606 76352 86674 76408
rect 86730 76352 86798 76408
rect 86854 76352 86922 76408
rect 86978 76352 87046 76408
rect 87102 76352 87126 76408
rect 86526 76284 87126 76352
rect 86526 76228 86550 76284
rect 86606 76228 86674 76284
rect 86730 76228 86798 76284
rect 86854 76228 86922 76284
rect 86978 76228 87046 76284
rect 87102 76228 87126 76284
rect 86526 76160 87126 76228
rect 86526 76104 86550 76160
rect 86606 76104 86674 76160
rect 86730 76104 86798 76160
rect 86854 76104 86922 76160
rect 86978 76104 87046 76160
rect 87102 76104 87126 76160
rect 86526 76036 87126 76104
rect 86526 75980 86550 76036
rect 86606 75980 86674 76036
rect 86730 75980 86798 76036
rect 86854 75980 86922 76036
rect 86978 75980 87046 76036
rect 87102 75980 87126 76036
rect 86526 75912 87126 75980
rect 86526 75856 86550 75912
rect 86606 75856 86674 75912
rect 86730 75856 86798 75912
rect 86854 75856 86922 75912
rect 86978 75856 87046 75912
rect 87102 75856 87126 75912
rect 86526 75788 87126 75856
rect 86526 75732 86550 75788
rect 86606 75732 86674 75788
rect 86730 75732 86798 75788
rect 86854 75732 86922 75788
rect 86978 75732 87046 75788
rect 87102 75732 87126 75788
rect 86526 63259 87126 75732
rect 86526 63203 86612 63259
rect 86668 63203 86736 63259
rect 86792 63203 86860 63259
rect 86916 63203 86984 63259
rect 87040 63203 87126 63259
rect 86526 63135 87126 63203
rect 86526 63079 86612 63135
rect 86668 63079 86736 63135
rect 86792 63079 86860 63135
rect 86916 63079 86984 63135
rect 87040 63079 87126 63135
rect 86526 63011 87126 63079
rect 86526 62955 86612 63011
rect 86668 62955 86736 63011
rect 86792 62955 86860 63011
rect 86916 62955 86984 63011
rect 87040 62955 87126 63011
rect 86526 62887 87126 62955
rect 86526 62831 86612 62887
rect 86668 62831 86736 62887
rect 86792 62831 86860 62887
rect 86916 62831 86984 62887
rect 87040 62831 87126 62887
rect 86526 61164 87126 62831
rect 86526 61108 86612 61164
rect 86668 61108 86736 61164
rect 86792 61108 86860 61164
rect 86916 61108 86984 61164
rect 87040 61108 87126 61164
rect 86526 61040 87126 61108
rect 86526 60984 86612 61040
rect 86668 60984 86736 61040
rect 86792 60984 86860 61040
rect 86916 60984 86984 61040
rect 87040 60984 87126 61040
rect 86526 60916 87126 60984
rect 86526 60860 86612 60916
rect 86668 60860 86736 60916
rect 86792 60860 86860 60916
rect 86916 60860 86984 60916
rect 87040 60860 87126 60916
rect 86526 60792 87126 60860
rect 86526 60736 86612 60792
rect 86668 60736 86736 60792
rect 86792 60736 86860 60792
rect 86916 60736 86984 60792
rect 87040 60736 87126 60792
rect 86526 59364 87126 60736
rect 86526 59308 86612 59364
rect 86668 59308 86736 59364
rect 86792 59308 86860 59364
rect 86916 59308 86984 59364
rect 87040 59308 87126 59364
rect 86526 59240 87126 59308
rect 86526 59184 86612 59240
rect 86668 59184 86736 59240
rect 86792 59184 86860 59240
rect 86916 59184 86984 59240
rect 87040 59184 87126 59240
rect 86526 59116 87126 59184
rect 86526 59060 86612 59116
rect 86668 59060 86736 59116
rect 86792 59060 86860 59116
rect 86916 59060 86984 59116
rect 87040 59060 87126 59116
rect 86526 58992 87126 59060
rect 86526 58936 86612 58992
rect 86668 58936 86736 58992
rect 86792 58936 86860 58992
rect 86916 58936 86984 58992
rect 87040 58936 87126 58992
rect 86526 57564 87126 58936
rect 86526 57508 86612 57564
rect 86668 57508 86736 57564
rect 86792 57508 86860 57564
rect 86916 57508 86984 57564
rect 87040 57508 87126 57564
rect 86526 57440 87126 57508
rect 86526 57384 86612 57440
rect 86668 57384 86736 57440
rect 86792 57384 86860 57440
rect 86916 57384 86984 57440
rect 87040 57384 87126 57440
rect 86526 57316 87126 57384
rect 86526 57260 86612 57316
rect 86668 57260 86736 57316
rect 86792 57260 86860 57316
rect 86916 57260 86984 57316
rect 87040 57260 87126 57316
rect 86526 57192 87126 57260
rect 86526 57136 86612 57192
rect 86668 57136 86736 57192
rect 86792 57136 86860 57192
rect 86916 57136 86984 57192
rect 87040 57136 87126 57192
rect 86526 55764 87126 57136
rect 86526 55708 86612 55764
rect 86668 55708 86736 55764
rect 86792 55708 86860 55764
rect 86916 55708 86984 55764
rect 87040 55708 87126 55764
rect 86526 55640 87126 55708
rect 86526 55584 86612 55640
rect 86668 55584 86736 55640
rect 86792 55584 86860 55640
rect 86916 55584 86984 55640
rect 87040 55584 87126 55640
rect 86526 55516 87126 55584
rect 86526 55460 86612 55516
rect 86668 55460 86736 55516
rect 86792 55460 86860 55516
rect 86916 55460 86984 55516
rect 87040 55460 87126 55516
rect 86526 55392 87126 55460
rect 86526 55336 86612 55392
rect 86668 55336 86736 55392
rect 86792 55336 86860 55392
rect 86916 55336 86984 55392
rect 87040 55336 87126 55392
rect 86526 53964 87126 55336
rect 86526 53908 86612 53964
rect 86668 53908 86736 53964
rect 86792 53908 86860 53964
rect 86916 53908 86984 53964
rect 87040 53908 87126 53964
rect 86526 53840 87126 53908
rect 86526 53784 86612 53840
rect 86668 53784 86736 53840
rect 86792 53784 86860 53840
rect 86916 53784 86984 53840
rect 87040 53784 87126 53840
rect 86526 53716 87126 53784
rect 86526 53660 86612 53716
rect 86668 53660 86736 53716
rect 86792 53660 86860 53716
rect 86916 53660 86984 53716
rect 87040 53660 87126 53716
rect 86526 53592 87126 53660
rect 86526 53536 86612 53592
rect 86668 53536 86736 53592
rect 86792 53536 86860 53592
rect 86916 53536 86984 53592
rect 87040 53536 87126 53592
rect 86526 52164 87126 53536
rect 86526 52108 86612 52164
rect 86668 52108 86736 52164
rect 86792 52108 86860 52164
rect 86916 52108 86984 52164
rect 87040 52108 87126 52164
rect 86526 52040 87126 52108
rect 86526 51984 86612 52040
rect 86668 51984 86736 52040
rect 86792 51984 86860 52040
rect 86916 51984 86984 52040
rect 87040 51984 87126 52040
rect 86526 51916 87126 51984
rect 86526 51860 86612 51916
rect 86668 51860 86736 51916
rect 86792 51860 86860 51916
rect 86916 51860 86984 51916
rect 87040 51860 87126 51916
rect 86526 51792 87126 51860
rect 86526 51736 86612 51792
rect 86668 51736 86736 51792
rect 86792 51736 86860 51792
rect 86916 51736 86984 51792
rect 87040 51736 87126 51792
rect 86526 50364 87126 51736
rect 86526 50308 86612 50364
rect 86668 50308 86736 50364
rect 86792 50308 86860 50364
rect 86916 50308 86984 50364
rect 87040 50308 87126 50364
rect 86526 50240 87126 50308
rect 86526 50184 86612 50240
rect 86668 50184 86736 50240
rect 86792 50184 86860 50240
rect 86916 50184 86984 50240
rect 87040 50184 87126 50240
rect 86526 50116 87126 50184
rect 86526 50060 86612 50116
rect 86668 50060 86736 50116
rect 86792 50060 86860 50116
rect 86916 50060 86984 50116
rect 87040 50060 87126 50116
rect 86526 49992 87126 50060
rect 86526 49936 86612 49992
rect 86668 49936 86736 49992
rect 86792 49936 86860 49992
rect 86916 49936 86984 49992
rect 87040 49936 87126 49992
rect 86526 48564 87126 49936
rect 86526 48508 86612 48564
rect 86668 48508 86736 48564
rect 86792 48508 86860 48564
rect 86916 48508 86984 48564
rect 87040 48508 87126 48564
rect 86526 48440 87126 48508
rect 86526 48384 86612 48440
rect 86668 48384 86736 48440
rect 86792 48384 86860 48440
rect 86916 48384 86984 48440
rect 87040 48384 87126 48440
rect 86526 48316 87126 48384
rect 86526 48260 86612 48316
rect 86668 48260 86736 48316
rect 86792 48260 86860 48316
rect 86916 48260 86984 48316
rect 87040 48260 87126 48316
rect 86526 48192 87126 48260
rect 86526 48136 86612 48192
rect 86668 48136 86736 48192
rect 86792 48136 86860 48192
rect 86916 48136 86984 48192
rect 87040 48136 87126 48192
rect 86526 46764 87126 48136
rect 86526 46708 86612 46764
rect 86668 46708 86736 46764
rect 86792 46708 86860 46764
rect 86916 46708 86984 46764
rect 87040 46708 87126 46764
rect 86526 46640 87126 46708
rect 86526 46584 86612 46640
rect 86668 46584 86736 46640
rect 86792 46584 86860 46640
rect 86916 46584 86984 46640
rect 87040 46584 87126 46640
rect 86526 46516 87126 46584
rect 86526 46460 86612 46516
rect 86668 46460 86736 46516
rect 86792 46460 86860 46516
rect 86916 46460 86984 46516
rect 87040 46460 87126 46516
rect 86526 46392 87126 46460
rect 86526 46336 86612 46392
rect 86668 46336 86736 46392
rect 86792 46336 86860 46392
rect 86916 46336 86984 46392
rect 87040 46336 87126 46392
rect 86526 44964 87126 46336
rect 86526 44908 86612 44964
rect 86668 44908 86736 44964
rect 86792 44908 86860 44964
rect 86916 44908 86984 44964
rect 87040 44908 87126 44964
rect 86526 44840 87126 44908
rect 86526 44784 86612 44840
rect 86668 44784 86736 44840
rect 86792 44784 86860 44840
rect 86916 44784 86984 44840
rect 87040 44784 87126 44840
rect 86526 44716 87126 44784
rect 86526 44660 86612 44716
rect 86668 44660 86736 44716
rect 86792 44660 86860 44716
rect 86916 44660 86984 44716
rect 87040 44660 87126 44716
rect 86526 44592 87126 44660
rect 86526 44536 86612 44592
rect 86668 44536 86736 44592
rect 86792 44536 86860 44592
rect 86916 44536 86984 44592
rect 87040 44536 87126 44592
rect 86526 43164 87126 44536
rect 86526 43108 86612 43164
rect 86668 43108 86736 43164
rect 86792 43108 86860 43164
rect 86916 43108 86984 43164
rect 87040 43108 87126 43164
rect 86526 43040 87126 43108
rect 86526 42984 86612 43040
rect 86668 42984 86736 43040
rect 86792 42984 86860 43040
rect 86916 42984 86984 43040
rect 87040 42984 87126 43040
rect 86526 42916 87126 42984
rect 86526 42860 86612 42916
rect 86668 42860 86736 42916
rect 86792 42860 86860 42916
rect 86916 42860 86984 42916
rect 87040 42860 87126 42916
rect 86526 42792 87126 42860
rect 86526 42736 86612 42792
rect 86668 42736 86736 42792
rect 86792 42736 86860 42792
rect 86916 42736 86984 42792
rect 87040 42736 87126 42792
rect 86526 41364 87126 42736
rect 86526 41308 86612 41364
rect 86668 41308 86736 41364
rect 86792 41308 86860 41364
rect 86916 41308 86984 41364
rect 87040 41308 87126 41364
rect 86526 41240 87126 41308
rect 86526 41184 86612 41240
rect 86668 41184 86736 41240
rect 86792 41184 86860 41240
rect 86916 41184 86984 41240
rect 87040 41184 87126 41240
rect 86526 41116 87126 41184
rect 86526 41060 86612 41116
rect 86668 41060 86736 41116
rect 86792 41060 86860 41116
rect 86916 41060 86984 41116
rect 87040 41060 87126 41116
rect 86526 40992 87126 41060
rect 86526 40936 86612 40992
rect 86668 40936 86736 40992
rect 86792 40936 86860 40992
rect 86916 40936 86984 40992
rect 87040 40936 87126 40992
rect 86526 39564 87126 40936
rect 86526 39508 86612 39564
rect 86668 39508 86736 39564
rect 86792 39508 86860 39564
rect 86916 39508 86984 39564
rect 87040 39508 87126 39564
rect 86526 39440 87126 39508
rect 86526 39384 86612 39440
rect 86668 39384 86736 39440
rect 86792 39384 86860 39440
rect 86916 39384 86984 39440
rect 87040 39384 87126 39440
rect 86526 39316 87126 39384
rect 86526 39260 86612 39316
rect 86668 39260 86736 39316
rect 86792 39260 86860 39316
rect 86916 39260 86984 39316
rect 87040 39260 87126 39316
rect 86526 39192 87126 39260
rect 86526 39136 86612 39192
rect 86668 39136 86736 39192
rect 86792 39136 86860 39192
rect 86916 39136 86984 39192
rect 87040 39136 87126 39192
rect 86526 37764 87126 39136
rect 86526 37708 86612 37764
rect 86668 37708 86736 37764
rect 86792 37708 86860 37764
rect 86916 37708 86984 37764
rect 87040 37708 87126 37764
rect 86526 37640 87126 37708
rect 86526 37584 86612 37640
rect 86668 37584 86736 37640
rect 86792 37584 86860 37640
rect 86916 37584 86984 37640
rect 87040 37584 87126 37640
rect 86526 37516 87126 37584
rect 86526 37460 86612 37516
rect 86668 37460 86736 37516
rect 86792 37460 86860 37516
rect 86916 37460 86984 37516
rect 87040 37460 87126 37516
rect 86526 37392 87126 37460
rect 86526 37336 86612 37392
rect 86668 37336 86736 37392
rect 86792 37336 86860 37392
rect 86916 37336 86984 37392
rect 87040 37336 87126 37392
rect 86526 35964 87126 37336
rect 86526 35908 86612 35964
rect 86668 35908 86736 35964
rect 86792 35908 86860 35964
rect 86916 35908 86984 35964
rect 87040 35908 87126 35964
rect 86526 35840 87126 35908
rect 86526 35784 86612 35840
rect 86668 35784 86736 35840
rect 86792 35784 86860 35840
rect 86916 35784 86984 35840
rect 87040 35784 87126 35840
rect 86526 35716 87126 35784
rect 86526 35660 86612 35716
rect 86668 35660 86736 35716
rect 86792 35660 86860 35716
rect 86916 35660 86984 35716
rect 87040 35660 87126 35716
rect 86526 35592 87126 35660
rect 86526 35536 86612 35592
rect 86668 35536 86736 35592
rect 86792 35536 86860 35592
rect 86916 35536 86984 35592
rect 87040 35536 87126 35592
rect 86526 34164 87126 35536
rect 86526 34108 86612 34164
rect 86668 34108 86736 34164
rect 86792 34108 86860 34164
rect 86916 34108 86984 34164
rect 87040 34108 87126 34164
rect 86526 34040 87126 34108
rect 86526 33984 86612 34040
rect 86668 33984 86736 34040
rect 86792 33984 86860 34040
rect 86916 33984 86984 34040
rect 87040 33984 87126 34040
rect 86526 33916 87126 33984
rect 86526 33860 86612 33916
rect 86668 33860 86736 33916
rect 86792 33860 86860 33916
rect 86916 33860 86984 33916
rect 87040 33860 87126 33916
rect 86526 33792 87126 33860
rect 86526 33736 86612 33792
rect 86668 33736 86736 33792
rect 86792 33736 86860 33792
rect 86916 33736 86984 33792
rect 87040 33736 87126 33792
rect 86526 32364 87126 33736
rect 86526 32308 86612 32364
rect 86668 32308 86736 32364
rect 86792 32308 86860 32364
rect 86916 32308 86984 32364
rect 87040 32308 87126 32364
rect 86526 32240 87126 32308
rect 86526 32184 86612 32240
rect 86668 32184 86736 32240
rect 86792 32184 86860 32240
rect 86916 32184 86984 32240
rect 87040 32184 87126 32240
rect 86526 32116 87126 32184
rect 86526 32060 86612 32116
rect 86668 32060 86736 32116
rect 86792 32060 86860 32116
rect 86916 32060 86984 32116
rect 87040 32060 87126 32116
rect 86526 31992 87126 32060
rect 86526 31936 86612 31992
rect 86668 31936 86736 31992
rect 86792 31936 86860 31992
rect 86916 31936 86984 31992
rect 87040 31936 87126 31992
rect 86526 30564 87126 31936
rect 86526 30508 86612 30564
rect 86668 30508 86736 30564
rect 86792 30508 86860 30564
rect 86916 30508 86984 30564
rect 87040 30508 87126 30564
rect 86526 30440 87126 30508
rect 86526 30384 86612 30440
rect 86668 30384 86736 30440
rect 86792 30384 86860 30440
rect 86916 30384 86984 30440
rect 87040 30384 87126 30440
rect 86526 30316 87126 30384
rect 86526 30260 86612 30316
rect 86668 30260 86736 30316
rect 86792 30260 86860 30316
rect 86916 30260 86984 30316
rect 87040 30260 87126 30316
rect 86526 30192 87126 30260
rect 86526 30136 86612 30192
rect 86668 30136 86736 30192
rect 86792 30136 86860 30192
rect 86916 30136 86984 30192
rect 87040 30136 87126 30192
rect 86526 28764 87126 30136
rect 86526 28708 86612 28764
rect 86668 28708 86736 28764
rect 86792 28708 86860 28764
rect 86916 28708 86984 28764
rect 87040 28708 87126 28764
rect 86526 28640 87126 28708
rect 86526 28584 86612 28640
rect 86668 28584 86736 28640
rect 86792 28584 86860 28640
rect 86916 28584 86984 28640
rect 87040 28584 87126 28640
rect 86526 28516 87126 28584
rect 86526 28460 86612 28516
rect 86668 28460 86736 28516
rect 86792 28460 86860 28516
rect 86916 28460 86984 28516
rect 87040 28460 87126 28516
rect 86526 28392 87126 28460
rect 86526 28336 86612 28392
rect 86668 28336 86736 28392
rect 86792 28336 86860 28392
rect 86916 28336 86984 28392
rect 87040 28336 87126 28392
rect 86526 26964 87126 28336
rect 86526 26908 86612 26964
rect 86668 26908 86736 26964
rect 86792 26908 86860 26964
rect 86916 26908 86984 26964
rect 87040 26908 87126 26964
rect 86526 26840 87126 26908
rect 86526 26784 86612 26840
rect 86668 26784 86736 26840
rect 86792 26784 86860 26840
rect 86916 26784 86984 26840
rect 87040 26784 87126 26840
rect 86526 26716 87126 26784
rect 86526 26660 86612 26716
rect 86668 26660 86736 26716
rect 86792 26660 86860 26716
rect 86916 26660 86984 26716
rect 87040 26660 87126 26716
rect 86526 26592 87126 26660
rect 86526 26536 86612 26592
rect 86668 26536 86736 26592
rect 86792 26536 86860 26592
rect 86916 26536 86984 26592
rect 87040 26536 87126 26592
rect 86526 25164 87126 26536
rect 86526 25108 86612 25164
rect 86668 25108 86736 25164
rect 86792 25108 86860 25164
rect 86916 25108 86984 25164
rect 87040 25108 87126 25164
rect 86526 25040 87126 25108
rect 86526 24984 86612 25040
rect 86668 24984 86736 25040
rect 86792 24984 86860 25040
rect 86916 24984 86984 25040
rect 87040 24984 87126 25040
rect 86526 24916 87126 24984
rect 86526 24860 86612 24916
rect 86668 24860 86736 24916
rect 86792 24860 86860 24916
rect 86916 24860 86984 24916
rect 87040 24860 87126 24916
rect 86526 24792 87126 24860
rect 86526 24736 86612 24792
rect 86668 24736 86736 24792
rect 86792 24736 86860 24792
rect 86916 24736 86984 24792
rect 87040 24736 87126 24792
rect 86526 23364 87126 24736
rect 86526 23308 86612 23364
rect 86668 23308 86736 23364
rect 86792 23308 86860 23364
rect 86916 23308 86984 23364
rect 87040 23308 87126 23364
rect 86526 23240 87126 23308
rect 86526 23184 86612 23240
rect 86668 23184 86736 23240
rect 86792 23184 86860 23240
rect 86916 23184 86984 23240
rect 87040 23184 87126 23240
rect 86526 23116 87126 23184
rect 86526 23060 86612 23116
rect 86668 23060 86736 23116
rect 86792 23060 86860 23116
rect 86916 23060 86984 23116
rect 87040 23060 87126 23116
rect 86526 22992 87126 23060
rect 86526 22936 86612 22992
rect 86668 22936 86736 22992
rect 86792 22936 86860 22992
rect 86916 22936 86984 22992
rect 87040 22936 87126 22992
rect 86526 21564 87126 22936
rect 86526 21508 86612 21564
rect 86668 21508 86736 21564
rect 86792 21508 86860 21564
rect 86916 21508 86984 21564
rect 87040 21508 87126 21564
rect 86526 21440 87126 21508
rect 86526 21384 86612 21440
rect 86668 21384 86736 21440
rect 86792 21384 86860 21440
rect 86916 21384 86984 21440
rect 87040 21384 87126 21440
rect 86526 21316 87126 21384
rect 86526 21260 86612 21316
rect 86668 21260 86736 21316
rect 86792 21260 86860 21316
rect 86916 21260 86984 21316
rect 87040 21260 87126 21316
rect 86526 21192 87126 21260
rect 86526 21136 86612 21192
rect 86668 21136 86736 21192
rect 86792 21136 86860 21192
rect 86916 21136 86984 21192
rect 87040 21136 87126 21192
rect 86526 19764 87126 21136
rect 86526 19708 86612 19764
rect 86668 19708 86736 19764
rect 86792 19708 86860 19764
rect 86916 19708 86984 19764
rect 87040 19708 87126 19764
rect 86526 19640 87126 19708
rect 86526 19584 86612 19640
rect 86668 19584 86736 19640
rect 86792 19584 86860 19640
rect 86916 19584 86984 19640
rect 87040 19584 87126 19640
rect 86526 19516 87126 19584
rect 86526 19460 86612 19516
rect 86668 19460 86736 19516
rect 86792 19460 86860 19516
rect 86916 19460 86984 19516
rect 87040 19460 87126 19516
rect 86526 19392 87126 19460
rect 86526 19336 86612 19392
rect 86668 19336 86736 19392
rect 86792 19336 86860 19392
rect 86916 19336 86984 19392
rect 87040 19336 87126 19392
rect 86526 17964 87126 19336
rect 86526 17908 86612 17964
rect 86668 17908 86736 17964
rect 86792 17908 86860 17964
rect 86916 17908 86984 17964
rect 87040 17908 87126 17964
rect 86526 17840 87126 17908
rect 86526 17784 86612 17840
rect 86668 17784 86736 17840
rect 86792 17784 86860 17840
rect 86916 17784 86984 17840
rect 87040 17784 87126 17840
rect 86526 17716 87126 17784
rect 86526 17660 86612 17716
rect 86668 17660 86736 17716
rect 86792 17660 86860 17716
rect 86916 17660 86984 17716
rect 87040 17660 87126 17716
rect 86526 17592 87126 17660
rect 86526 17536 86612 17592
rect 86668 17536 86736 17592
rect 86792 17536 86860 17592
rect 86916 17536 86984 17592
rect 87040 17536 87126 17592
rect 86526 16164 87126 17536
rect 86526 16108 86612 16164
rect 86668 16108 86736 16164
rect 86792 16108 86860 16164
rect 86916 16108 86984 16164
rect 87040 16108 87126 16164
rect 86526 16040 87126 16108
rect 86526 15984 86612 16040
rect 86668 15984 86736 16040
rect 86792 15984 86860 16040
rect 86916 15984 86984 16040
rect 87040 15984 87126 16040
rect 86526 15916 87126 15984
rect 86526 15860 86612 15916
rect 86668 15860 86736 15916
rect 86792 15860 86860 15916
rect 86916 15860 86984 15916
rect 87040 15860 87126 15916
rect 86526 15792 87126 15860
rect 86526 15736 86612 15792
rect 86668 15736 86736 15792
rect 86792 15736 86860 15792
rect 86916 15736 86984 15792
rect 87040 15736 87126 15792
rect 86526 14364 87126 15736
rect 86526 14308 86612 14364
rect 86668 14308 86736 14364
rect 86792 14308 86860 14364
rect 86916 14308 86984 14364
rect 87040 14308 87126 14364
rect 86526 14240 87126 14308
rect 86526 14184 86612 14240
rect 86668 14184 86736 14240
rect 86792 14184 86860 14240
rect 86916 14184 86984 14240
rect 87040 14184 87126 14240
rect 86526 14116 87126 14184
rect 86526 14060 86612 14116
rect 86668 14060 86736 14116
rect 86792 14060 86860 14116
rect 86916 14060 86984 14116
rect 87040 14060 87126 14116
rect 86526 13992 87126 14060
rect 86526 13936 86612 13992
rect 86668 13936 86736 13992
rect 86792 13936 86860 13992
rect 86916 13936 86984 13992
rect 87040 13936 87126 13992
rect 86526 12564 87126 13936
rect 86526 12508 86612 12564
rect 86668 12508 86736 12564
rect 86792 12508 86860 12564
rect 86916 12508 86984 12564
rect 87040 12508 87126 12564
rect 86526 12440 87126 12508
rect 86526 12384 86612 12440
rect 86668 12384 86736 12440
rect 86792 12384 86860 12440
rect 86916 12384 86984 12440
rect 87040 12384 87126 12440
rect 86526 12316 87126 12384
rect 86526 12260 86612 12316
rect 86668 12260 86736 12316
rect 86792 12260 86860 12316
rect 86916 12260 86984 12316
rect 87040 12260 87126 12316
rect 86526 12192 87126 12260
rect 86526 12136 86612 12192
rect 86668 12136 86736 12192
rect 86792 12136 86860 12192
rect 86916 12136 86984 12192
rect 87040 12136 87126 12192
rect 86526 10764 87126 12136
rect 86526 10708 86612 10764
rect 86668 10708 86736 10764
rect 86792 10708 86860 10764
rect 86916 10708 86984 10764
rect 87040 10708 87126 10764
rect 86526 10640 87126 10708
rect 86526 10584 86612 10640
rect 86668 10584 86736 10640
rect 86792 10584 86860 10640
rect 86916 10584 86984 10640
rect 87040 10584 87126 10640
rect 86526 10516 87126 10584
rect 86526 10460 86612 10516
rect 86668 10460 86736 10516
rect 86792 10460 86860 10516
rect 86916 10460 86984 10516
rect 87040 10460 87126 10516
rect 86526 10392 87126 10460
rect 86526 10336 86612 10392
rect 86668 10336 86736 10392
rect 86792 10336 86860 10392
rect 86916 10336 86984 10392
rect 87040 10336 87126 10392
rect 86526 8964 87126 10336
rect 86526 8908 86612 8964
rect 86668 8908 86736 8964
rect 86792 8908 86860 8964
rect 86916 8908 86984 8964
rect 87040 8908 87126 8964
rect 86526 8840 87126 8908
rect 86526 8784 86612 8840
rect 86668 8784 86736 8840
rect 86792 8784 86860 8840
rect 86916 8784 86984 8840
rect 87040 8784 87126 8840
rect 86526 8716 87126 8784
rect 86526 8660 86612 8716
rect 86668 8660 86736 8716
rect 86792 8660 86860 8716
rect 86916 8660 86984 8716
rect 87040 8660 87126 8716
rect 86526 8592 87126 8660
rect 86526 8536 86612 8592
rect 86668 8536 86736 8592
rect 86792 8536 86860 8592
rect 86916 8536 86984 8592
rect 87040 8536 87126 8592
rect 86526 7164 87126 8536
rect 86526 7108 86612 7164
rect 86668 7108 86736 7164
rect 86792 7108 86860 7164
rect 86916 7108 86984 7164
rect 87040 7108 87126 7164
rect 86526 7040 87126 7108
rect 86526 6984 86612 7040
rect 86668 6984 86736 7040
rect 86792 6984 86860 7040
rect 86916 6984 86984 7040
rect 87040 6984 87126 7040
rect 86526 6916 87126 6984
rect 86526 6860 86612 6916
rect 86668 6860 86736 6916
rect 86792 6860 86860 6916
rect 86916 6860 86984 6916
rect 87040 6860 87126 6916
rect 86526 6792 87126 6860
rect 86526 6736 86612 6792
rect 86668 6736 86736 6792
rect 86792 6736 86860 6792
rect 86916 6736 86984 6792
rect 87040 6736 87126 6792
rect 86526 5364 87126 6736
rect 86526 5308 86612 5364
rect 86668 5308 86736 5364
rect 86792 5308 86860 5364
rect 86916 5308 86984 5364
rect 87040 5308 87126 5364
rect 86526 5240 87126 5308
rect 86526 5184 86612 5240
rect 86668 5184 86736 5240
rect 86792 5184 86860 5240
rect 86916 5184 86984 5240
rect 87040 5184 87126 5240
rect 86526 5116 87126 5184
rect 86526 5060 86612 5116
rect 86668 5060 86736 5116
rect 86792 5060 86860 5116
rect 86916 5060 86984 5116
rect 87040 5060 87126 5116
rect 86526 4992 87126 5060
rect 86526 4936 86612 4992
rect 86668 4936 86736 4992
rect 86792 4936 86860 4992
rect 86916 4936 86984 4992
rect 87040 4936 87126 4992
rect 86526 3632 87126 4936
rect 86526 3576 86612 3632
rect 86668 3576 86736 3632
rect 86792 3576 86860 3632
rect 86916 3576 86984 3632
rect 87040 3576 87126 3632
rect 86526 3508 87126 3576
rect 86526 3452 86612 3508
rect 86668 3452 86736 3508
rect 86792 3452 86860 3508
rect 86916 3452 86984 3508
rect 87040 3452 87126 3508
rect 86526 3384 87126 3452
rect 86526 3328 86612 3384
rect 86668 3328 86736 3384
rect 86792 3328 86860 3384
rect 86916 3328 86984 3384
rect 87040 3328 87126 3384
rect 86526 3260 87126 3328
rect 86526 3204 86612 3260
rect 86668 3204 86736 3260
rect 86792 3204 86860 3260
rect 86916 3204 86984 3260
rect 87040 3204 87126 3260
rect 86526 3136 87126 3204
use gf180mcu_fd_ip_sram__sram512x8m8wm1  sram512x8
timestamp 0
transform -1 0 87372 0 -1 97976
box 0 0 86372 96976
<< labels >>
flabel metal2 s 52944 98376 53056 99176 0 FreeSans 448 90 0 0 A[0]
port 0 nsew signal input
flabel metal2 s 54644 98376 54756 99176 0 FreeSans 448 90 0 0 A[1]
port 1 nsew signal input
flabel metal2 s 56344 98376 56456 99176 0 FreeSans 448 90 0 0 A[2]
port 2 nsew signal input
flabel metal2 s 30944 98376 31056 99176 0 FreeSans 448 90 0 0 A[3]
port 3 nsew signal input
flabel metal2 s 31944 98376 32056 99176 0 FreeSans 448 90 0 0 A[4]
port 4 nsew signal input
flabel metal2 s 32744 98376 32856 99176 0 FreeSans 448 90 0 0 A[5]
port 5 nsew signal input
flabel metal2 s 33344 98376 33456 99176 0 FreeSans 448 90 0 0 A[6]
port 6 nsew signal input
flabel metal2 s 57444 98376 57556 99176 0 FreeSans 448 90 0 0 A[7]
port 7 nsew signal input
flabel metal2 s 58144 98376 58256 99176 0 FreeSans 448 90 0 0 A[8]
port 8 nsew signal input
flabel metal2 s 36844 98376 36956 99176 0 FreeSans 448 90 0 0 CEN
port 9 nsew signal input
flabel metal2 s 59244 98376 59356 99176 0 FreeSans 448 90 0 0 CLK
port 10 nsew signal input
flabel metal2 s 85344 98376 85456 99176 0 FreeSans 448 90 0 0 D[0]
port 11 nsew signal input
flabel metal2 s 74944 98376 75056 99176 0 FreeSans 448 90 0 0 D[1]
port 12 nsew signal input
flabel metal2 s 73744 98376 73856 99176 0 FreeSans 448 90 0 0 D[2]
port 13 nsew signal input
flabel metal2 s 63344 98376 63456 99176 0 FreeSans 448 90 0 0 D[3]
port 14 nsew signal input
flabel metal2 s 25744 98376 25856 99176 0 FreeSans 448 90 0 0 D[4]
port 15 nsew signal input
flabel metal2 s 15444 98376 15556 99176 0 FreeSans 448 90 0 0 D[5]
port 16 nsew signal input
flabel metal2 s 14144 98376 14256 99176 0 FreeSans 448 90 0 0 D[6]
port 17 nsew signal input
flabel metal2 s 3744 98376 3856 99176 0 FreeSans 448 90 0 0 D[7]
port 18 nsew signal input
flabel metal2 s 46568 98376 46680 99176 0 FreeSans 448 90 0 0 GWEN
port 19 nsew signal input
flabel metal2 s 83844 98376 83956 99176 0 FreeSans 448 90 0 0 Q[0]
port 20 nsew signal tristate
flabel metal2 s 75644 98376 75756 99176 0 FreeSans 448 90 0 0 Q[1]
port 21 nsew signal tristate
flabel metal2 s 73044 98376 73156 99176 0 FreeSans 448 90 0 0 Q[2]
port 22 nsew signal tristate
flabel metal2 s 64944 98376 65056 99176 0 FreeSans 448 90 0 0 Q[3]
port 23 nsew signal tristate
flabel metal2 s 24244 98376 24356 99176 0 FreeSans 448 90 0 0 Q[4]
port 24 nsew signal tristate
flabel metal2 s 16044 98376 16156 99176 0 FreeSans 448 90 0 0 Q[5]
port 25 nsew signal tristate
flabel metal2 s 13444 98376 13556 99176 0 FreeSans 448 90 0 0 Q[6]
port 26 nsew signal tristate
flabel metal2 s 5344 98376 5456 99176 0 FreeSans 448 90 0 0 Q[7]
port 27 nsew signal tristate
flabel metal4 s 1044 3136 1644 95648 0 FreeSans 2560 90 0 0 VDD
port 28 nsew power bidirectional
flabel metal4 s 85726 3136 86326 95648 0 FreeSans 2560 90 0 0 VDD
port 28 nsew power bidirectional
flabel metal4 s 1844 3136 2444 95648 0 FreeSans 2560 90 0 0 VSS
port 29 nsew ground bidirectional
flabel metal4 s 86526 3136 87126 95648 0 FreeSans 2560 90 0 0 VSS
port 29 nsew ground bidirectional
flabel metal2 s 84644 98376 84756 99176 0 FreeSans 448 90 0 0 WEN[0]
port 30 nsew signal input
flabel metal2 s 74544 98376 74656 99176 0 FreeSans 448 90 0 0 WEN[1]
port 31 nsew signal input
flabel metal2 s 74144 98376 74256 99176 0 FreeSans 448 90 0 0 WEN[2]
port 32 nsew signal input
flabel metal2 s 63744 98376 63856 99176 0 FreeSans 448 90 0 0 WEN[3]
port 33 nsew signal input
flabel metal2 s 25044 98376 25156 99176 0 FreeSans 448 90 0 0 WEN[4]
port 34 nsew signal input
flabel metal2 s 14994 98376 15106 99176 0 FreeSans 448 90 0 0 WEN[5]
port 35 nsew signal input
flabel metal2 s 14544 98376 14656 99176 0 FreeSans 448 90 0 0 WEN[6]
port 36 nsew signal input
flabel metal2 s 4444 98376 4556 99176 0 FreeSans 448 90 0 0 WEN[7]
port 37 nsew signal input
rlabel via3 86274 89763 86274 89763 0 VDD
rlabel via3 87074 95397 87074 95397 0 VSS
rlabel metal2 53032 98224 53032 98224 0 A[0]
rlabel metal2 54712 98224 54712 98224 0 A[1]
rlabel metal2 56392 98224 56392 98224 0 A[2]
rlabel metal2 30968 98224 30968 98224 0 A[3]
rlabel metal2 32032 98070 32032 98070 0 A[4]
rlabel metal2 32760 98224 32760 98224 0 A[5]
rlabel metal2 33432 98224 33432 98224 0 A[6]
rlabel metal2 57512 98224 57512 98224 0 A[7]
rlabel metal2 58184 98224 58184 98224 0 A[8]
rlabel metal2 36904 98224 36904 98224 0 CEN
rlabel metal2 59304 98224 59304 98224 0 CLK
rlabel metal2 85400 98224 85400 98224 0 D[0]
rlabel metal2 74984 98224 74984 98224 0 D[1]
rlabel metal2 73752 98224 73752 98224 0 D[2]
rlabel metal2 63448 98224 63448 98224 0 D[3]
rlabel metal2 25816 98224 25816 98224 0 D[4]
rlabel metal2 15512 98224 15512 98224 0 D[5]
rlabel metal2 14168 98224 14168 98224 0 D[6]
rlabel metal2 3808 98070 3808 98070 0 D[7]
rlabel metal2 46648 98224 46648 98224 0 GWEN
rlabel metal2 83944 98224 83944 98224 0 Q[0]
rlabel metal2 75656 98224 75656 98224 0 Q[1]
rlabel metal2 73080 98224 73080 98224 0 Q[2]
rlabel metal2 65016 98224 65016 98224 0 Q[3]
rlabel metal2 24248 98224 24248 98224 0 Q[4]
rlabel metal2 16072 98224 16072 98224 0 Q[5]
rlabel metal2 13496 98224 13496 98224 0 Q[6]
rlabel metal2 5432 98224 5432 98224 0 Q[7]
rlabel metal2 84728 98224 84728 98224 0 WEN[0]
rlabel metal2 74648 98224 74648 98224 0 WEN[1]
rlabel metal2 74200 98224 74200 98224 0 WEN[2]
rlabel metal2 63784 98224 63784 98224 0 WEN[3]
rlabel metal2 25144 98224 25144 98224 0 WEN[4]
rlabel metal2 15064 98224 15064 98224 0 WEN[5]
rlabel metal2 14616 98224 14616 98224 0 WEN[6]
rlabel metal2 4536 98224 4536 98224 0 WEN[7]
<< properties >>
string FIXED_BBOX 0 0 88972 99176
<< end >>
