// This is the unpowered netlist.
module gpios (DAC_clk,
    DAC_d1,
    DAC_d2,
    DAC_le,
    RXD,
    TXD,
    bus_cyc,
    bus_we,
    irq0,
    irq6,
    irq7,
    pwm0,
    pwm1,
    pwm2,
    rst,
    tmr0_clk,
    tmr0_o,
    tmr1_clk,
    tmr1_o,
    wb_clk_i,
    addr,
    data_in,
    data_out,
    io_in,
    io_oeb,
    io_out,
    la_data_out);
 input DAC_clk;
 input DAC_d1;
 input DAC_d2;
 input DAC_le;
 output RXD;
 input TXD;
 input bus_cyc;
 input bus_we;
 output irq0;
 output irq6;
 output irq7;
 input pwm0;
 input pwm1;
 input pwm2;
 input rst;
 output tmr0_clk;
 input tmr0_o;
 output tmr1_clk;
 input tmr1_o;
 input wb_clk_i;
 input [3:0] addr;
 input [7:0] data_in;
 output [7:0] data_out;
 input [15:0] io_in;
 output [15:0] io_oeb;
 output [15:0] io_out;
 output [7:0] la_data_out;

 wire \DDRA[0] ;
 wire \DDRA[1] ;
 wire \DDRA[2] ;
 wire \DDRA[3] ;
 wire \DDRA[4] ;
 wire \DDRA[5] ;
 wire \DDRA[6] ;
 wire \DDRA[7] ;
 wire \DDRB[0] ;
 wire \DDRB[1] ;
 wire \DDRB[2] ;
 wire \DDRB[3] ;
 wire \DDRB[4] ;
 wire \DDRB[5] ;
 wire \DDRB[6] ;
 wire \DDRB[7] ;
 wire \PORTA[0] ;
 wire \PORTA[1] ;
 wire \PORTA[2] ;
 wire \PORTA[3] ;
 wire \PORTA[4] ;
 wire \PORTA[5] ;
 wire \PORTA[6] ;
 wire \PORTA[7] ;
 wire \PORTB[0] ;
 wire \PORTB[1] ;
 wire \PORTB[2] ;
 wire \PORTB[3] ;
 wire \PORTB[4] ;
 wire \PORTB[5] ;
 wire \PORTB[6] ;
 wire \PORTB[7] ;
 wire \SPA[0] ;
 wire \SPA[1] ;
 wire \SPA[2] ;
 wire \SPA[3] ;
 wire \SPA[4] ;
 wire \SPA[5] ;
 wire \SPA[6] ;
 wire \SPA[7] ;
 wire \SPB[0] ;
 wire \SPB[1] ;
 wire \SPB[2] ;
 wire \SPB[3] ;
 wire \SPB[4] ;
 wire \SPB[5] ;
 wire \SPB[6] ;
 wire \SPB[7] ;
 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire _172_;
 wire _173_;
 wire _174_;
 wire _175_;
 wire _176_;
 wire _177_;
 wire _178_;
 wire _179_;
 wire _180_;
 wire _181_;
 wire _182_;
 wire _183_;
 wire _184_;
 wire _185_;
 wire _186_;
 wire _187_;
 wire _188_;
 wire _189_;
 wire _190_;
 wire _191_;
 wire _192_;
 wire _193_;
 wire _194_;
 wire _195_;
 wire _196_;
 wire _197_;
 wire _198_;
 wire _199_;
 wire _200_;
 wire _201_;
 wire _202_;
 wire _203_;
 wire _204_;
 wire _205_;
 wire _206_;
 wire _207_;
 wire _208_;
 wire _209_;
 wire _210_;
 wire _211_;
 wire _212_;
 wire _213_;
 wire _214_;
 wire _215_;
 wire _216_;
 wire _217_;
 wire _218_;
 wire _219_;
 wire _220_;
 wire _221_;
 wire _222_;
 wire _223_;
 wire _224_;
 wire _225_;
 wire _226_;
 wire _227_;
 wire _228_;
 wire _229_;
 wire _230_;
 wire _231_;
 wire _232_;
 wire _233_;
 wire _234_;
 wire _235_;
 wire _236_;
 wire _237_;
 wire _238_;
 wire _239_;
 wire _240_;
 wire _241_;
 wire _242_;
 wire _243_;
 wire _244_;
 wire _245_;
 wire _246_;
 wire _247_;
 wire _248_;
 wire _249_;
 wire _250_;
 wire _251_;
 wire _252_;
 wire _253_;
 wire _254_;
 wire _255_;
 wire _256_;
 wire _257_;
 wire _258_;
 wire _259_;
 wire _260_;
 wire _261_;
 wire _262_;
 wire _263_;
 wire _264_;
 wire _265_;
 wire _266_;
 wire _267_;
 wire _268_;
 wire _269_;
 wire _270_;
 wire _271_;
 wire _272_;
 wire _273_;
 wire _274_;
 wire _275_;
 wire _276_;
 wire _277_;
 wire _278_;
 wire _279_;
 wire _280_;
 wire _281_;
 wire _282_;
 wire _283_;
 wire _284_;
 wire _285_;
 wire _286_;
 wire _287_;
 wire _288_;
 wire _289_;
 wire _290_;
 wire _291_;
 wire _292_;
 wire _293_;
 wire _294_;
 wire _295_;
 wire _296_;
 wire _297_;
 wire _298_;
 wire _299_;
 wire _300_;
 wire _301_;
 wire _302_;
 wire _303_;
 wire _304_;
 wire _305_;
 wire _306_;
 wire _307_;
 wire _308_;
 wire _309_;
 wire _310_;
 wire _311_;
 wire _312_;
 wire _313_;
 wire _314_;
 wire _315_;
 wire _316_;
 wire _317_;
 wire _318_;
 wire _319_;
 wire _320_;
 wire _321_;
 wire _322_;
 wire _323_;
 wire _324_;
 wire _325_;
 wire _326_;
 wire _327_;
 wire _328_;
 wire _329_;
 wire _330_;
 wire _331_;
 wire _332_;
 wire _333_;
 wire _334_;
 wire _335_;
 wire _336_;
 wire _337_;
 wire _338_;
 wire _339_;
 wire _340_;
 wire _341_;
 wire _342_;
 wire _343_;
 wire _344_;
 wire _345_;
 wire _346_;
 wire _347_;
 wire _348_;
 wire _349_;
 wire _350_;
 wire _351_;
 wire _352_;
 wire _353_;
 wire _354_;
 wire _355_;
 wire _356_;
 wire _357_;
 wire _358_;
 wire _359_;
 wire _360_;
 wire _361_;
 wire _362_;
 wire _363_;
 wire _364_;
 wire _365_;
 wire _366_;
 wire _367_;
 wire _368_;
 wire _369_;
 wire _370_;
 wire _371_;
 wire _372_;
 wire _373_;
 wire _374_;
 wire _375_;
 wire _376_;
 wire _377_;
 wire _378_;
 wire _379_;
 wire _380_;
 wire _381_;
 wire _382_;
 wire _383_;
 wire _384_;
 wire _385_;
 wire _386_;
 wire _387_;
 wire _388_;
 wire _389_;
 wire _390_;
 wire _391_;
 wire _392_;
 wire _393_;
 wire _394_;
 wire _395_;
 wire _396_;
 wire _397_;
 wire _398_;
 wire _399_;
 wire clknet_0_wb_clk_i;
 wire clknet_3_0__leaf_wb_clk_i;
 wire clknet_3_1__leaf_wb_clk_i;
 wire clknet_3_2__leaf_wb_clk_i;
 wire clknet_3_3__leaf_wb_clk_i;
 wire clknet_3_4__leaf_wb_clk_i;
 wire clknet_3_5__leaf_wb_clk_i;
 wire clknet_3_6__leaf_wb_clk_i;
 wire clknet_3_7__leaf_wb_clk_i;
 wire last_irg6_trigger;
 wire last_irq0_trigger;
 wire last_irq7_trigger;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;

 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__401__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__I1 (.I(net5));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__403__S (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__405__I (.I(\SPA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__406__A2 (.I(\PORTA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__I0 (.I(\PORTA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__I1 (.I(net40));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__408__S (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__I0 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__I1 (.I(net41));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__410__S (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__I0 (.I(\PORTA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__I1 (.I(net36));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__412__S (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__I0 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__I1 (.I(net37));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__414__S (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__416__I (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__419__A1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__420__A2 (.I(\DDRA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__421__A2 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__A1 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__422__A2 (.I(\DDRA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__423__A2 (.I(\DDRA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__A1 (.I(\SPA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__425__A2 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__429__S (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__433__A2 (.I(_086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__434__I (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__435__A2 (.I(\PORTB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__I0 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__437__S (.I(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__I0 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__439__S (.I(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__I0 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__441__S (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__I0 (.I(\PORTB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__443__S (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A1 (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__445__A2 (.I(\DDRB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__446__A1 (.I(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A1 (.I(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__447__A2 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A1 (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__448__A2 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A1 (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__449__A2 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__450__A2 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__451__A2 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__453__A2 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__455__A2 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__457__A2 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__458__A2 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__460__A1 (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__461__I (.I(_096_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__462__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__464__I (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A1 (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__465__A2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__466__A2 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__467__I (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__468__I (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__472__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__473__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__474__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__475__A3 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__477__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__478__I (.I(net6));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__480__I (.I(net7));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__482__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__484__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__B2 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__490__C2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__491__A1 (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__494__I (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A1 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__495__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__496__I (.I(net8));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__497__I (.I(net9));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__502__I (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__504__I (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A1 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__A2 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__511__B2 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__514__C (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A1 (.I(\DDRB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__517__A2 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__A2 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__519__C1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__521__I (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__522__I (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__523__A1 (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__525__C (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__529__B2 (.I(_081_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__531__I (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__533__I (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__A1 (.I(net21));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__534__C1 (.I(\SPA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__535__I (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__A1 (.I(\PORTA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__A2 (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__536__B2 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__542__I (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__A1 (.I(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__B2 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__544__C2 (.I(\DDRA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__A2 (.I(_140_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__B1 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__B2 (.I(\PORTA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__545__C1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__546__A1 (.I(\PORTB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__A1 (.I(_181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__553__B2 (.I(_182_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__A1 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__554__B2 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__B1 (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__B2 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__555__C1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__556__A1 (.I(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__A1 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__B2 (.I(\DDRA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__560__C2 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__561__A1 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A1 (.I(\PORTA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__A2 (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__562__B2 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__563__A1 (.I(net24));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__A1 (.I(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__564__B2 (.I(net31));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__A1 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__B2 (.I(\DDRA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__568__C2 (.I(net32));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__B2 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__569__C1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__570__A1 (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__571__A1 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__571__B2 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__573__C (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__577__C (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__A1 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__578__B2 (.I(net33));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__579__B2 (.I(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__580__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__A1 (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__B2 (.I(\PORTB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__581__C1 (.I(_167_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__583__C (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__584__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A1 (.I(net10));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__585__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A1 (.I(_210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__588__A3 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__589__A2 (.I(net20));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__591__A1 (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__593__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A1 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__594__A3 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__595__A2 (.I(net34));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__597__A1 (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__599__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__600__A3 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__601__A2 (.I(_100_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__602__A1 (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__604__I (.I(net12));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__606__A1 (.I(_101_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__606__A2 (.I(net11));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__609__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__611__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__615__I (.I(_098_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__618__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__620__C (.I(_241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__621__I (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__622__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__627__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__628__C (.I(_241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__629__I (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__630__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__634__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__635__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__637__C (.I(_254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__638__I (.I(net18));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__639__A1 (.I(_255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__642__I (.I(net19));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__643__A1 (.I(_258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__645__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__647__B (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__649__A2 (.I(_263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__651__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__652__A2 (.I(_213_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__654__A1 (.I(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__655__B (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__656__I (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__657__A1 (.I(_270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__659__B (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__660__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__661__A1 (.I(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__662__B (.I(_262_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__663__I (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__664__A1 (.I(_275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__665__A1 (.I(\DDRA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__669__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__671__A1 (.I(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__673__I (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__674__A1 (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__675__A1 (.I(\DDRA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__677__A1 (.I(_255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__678__A1 (.I(\DDRA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__680__A1 (.I(_258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__686__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__687__A1 (.I(_126_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__690__A1 (.I(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__692__I (.I(\DDRB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__693__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__694__C (.I(_254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__695__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__696__A1 (.I(_093_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__696__C (.I(_254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__697__A1 (.I(_275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__699__A1 (.I(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__701__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__702__A1 (.I(_181_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__702__C (.I(_254_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__703__A1 (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__704__A1 (.I(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__706__A1 (.I(_255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__707__A1 (.I(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__709__B (.I(_309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__710__A1 (.I(_258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__711__A1 (.I(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__712__B (.I(_309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__A1 (.I(_135_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__713__A2 (.I(_263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__715__A1 (.I(_227_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__716__A2 (.I(_263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__719__B (.I(_309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__720__A1 (.I(_270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__722__B (.I(_309_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__723__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__724__A1 (.I(\PORTA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__725__I (.I(net39));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__728__A1 (.I(_275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__729__A1 (.I(\PORTA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__732__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__734__A1 (.I(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__736__A1 (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__737__A1 (.I(\PORTA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__739__A1 (.I(_255_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__740__A1 (.I(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__743__A1 (.I(_258_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__746__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__748__A1 (.I(_210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__749__A1 (.I(_127_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__753__A1 (.I(_270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__756__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__758__A1 (.I(_086_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__759__A1 (.I(_275_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__760__A1 (.I(\PORTB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__763__A1 (.I(_248_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__765__A1 (.I(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__767__A1 (.I(_283_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__768__A1 (.I(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__770__A1 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__771__A1 (.I(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__773__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__774__A1 (.I(\PORTB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__776__B (.I(_359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__777__A1 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__780__A1 (.I(_210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__781__A1 (.I(_070_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__782__A1 (.I(_137_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__782__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__784__A1 (.I(_270_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__785__A1 (.I(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__786__B (.I(_359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__787__A1 (.I(net14));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__788__A1 (.I(_073_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__789__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__791__A1 (.I(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__792__B (.I(_359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__793__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__794__A1 (.I(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__795__B (.I(_359_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__796__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__797__A1 (.I(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__800__A1 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__801__A1 (.I(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__803__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__805__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__805__A2 (.I(_263_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__807__A1 (.I(_210_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__808__C (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__809__A1 (.I(_110_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__809__A2 (.I(_233_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__811__A1 (.I(net13));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__812__A1 (.I(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__814__A1 (.I(_242_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__815__A1 (.I(_085_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__817__A1 (.I(net15));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__818__C (.I(_147_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__819__A1 (.I(net16));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__821__A1 (.I(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__824__A1 (.I(net17));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__825__A1 (.I(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__827__A1 (.I(_218_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__828__A1 (.I(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__830__A1 (.I(_223_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__831__A1 (.I(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__833__A1 (.I(_241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__834__A1 (.I(_241_));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__835__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__836__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__837__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__838__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__839__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__840__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__841__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__842__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__843__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__844__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__845__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__846__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__847__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__848__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__849__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__850__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__851__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__852__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__853__CLK (.I(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__854__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__855__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__856__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__857__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__858__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__859__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__860__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__861__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__862__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__863__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__864__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__865__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__866__CLK (.I(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__867__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__868__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__869__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__870__CLK (.I(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__871__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__872__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__873__CLK (.I(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__874__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__875__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__876__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__877__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__878__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__879__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__880__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__881__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__882__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__883__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__884__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__885__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__886__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__887__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__888__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__889__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__890__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__891__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__892__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__893__CLK (.I(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__894__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__895__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__896__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__897__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__898__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__899__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__900__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__901__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__902__CLK (.I(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__903__CLK (.I(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA__904__CLK (.I(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_0_wb_clk_i_I (.I(wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_0__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_1__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_2__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_3__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_4__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_5__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_6__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_clkbuf_3_7__f_wb_clk_i_I (.I(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input10_I (.I(bus_cyc));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input11_I (.I(bus_we));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input12_I (.I(data_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input13_I (.I(data_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input14_I (.I(data_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input15_I (.I(data_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input16_I (.I(data_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input17_I (.I(data_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input18_I (.I(data_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input19_I (.I(data_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input1_I (.I(DAC_clk));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input20_I (.I(io_in[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input21_I (.I(io_in[10]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input22_I (.I(io_in[11]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input23_I (.I(io_in[12]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input24_I (.I(io_in[13]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input25_I (.I(io_in[14]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input26_I (.I(io_in[15]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input27_I (.I(io_in[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input28_I (.I(io_in[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input29_I (.I(io_in[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input2_I (.I(DAC_d1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input30_I (.I(io_in[4]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input31_I (.I(io_in[5]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input32_I (.I(io_in[6]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input33_I (.I(io_in[7]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input34_I (.I(io_in[8]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input35_I (.I(io_in[9]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input36_I (.I(pwm0));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input37_I (.I(pwm1));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input38_I (.I(pwm2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input39_I (.I(rst));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input3_I (.I(DAC_d2));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input40_I (.I(tmr0_o));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input41_I (.I(tmr1_o));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input4_I (.I(DAC_le));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input5_I (.I(TXD));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input6_I (.I(addr[0]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input7_I (.I(addr[1]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input8_I (.I(addr[2]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_input9_I (.I(addr[3]));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output53_I (.I(net53));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output64_I (.I(net64));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output65_I (.I(net65));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output83_I (.I(net83));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output84_I (.I(net84));
 gf180mcu_fd_sc_mcu7t5v0__antenna ANTENNA_output85_I (.I(net85));
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_0_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_0_339 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_418 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_0_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_0_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_10_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_10_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_10_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_10_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_10_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_10_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_10_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_11_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_11_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_11_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_11_38 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_11_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_11_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_11_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_12_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_12_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_12_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_12_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_12_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_12_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_12_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_13_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_13_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_13_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_13_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_13_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_13_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_13_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_14_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_14_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_14_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_14_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_14_75 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_14_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_14_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_15_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_15_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_15_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_15_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_15_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_15_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_16_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_16_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_16_71 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_16_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_16_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_16_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_14 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_159 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_318 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_17_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_17_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_17_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_17_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_17_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_17_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_17_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_213 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_18_275 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_18_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_18_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_18_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_18_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_18_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_18_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_19_332 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_19_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_50 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_19_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_19_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_19_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_19_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_24 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_1_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_354 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_1_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_397 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_405 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_1_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_1_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_1_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_1_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_322 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_326 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_330 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_20_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_378 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_20_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_20_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_20_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_20_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_20_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_269 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_21_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_21_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_21_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_21_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_21_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_21_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_109 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_302 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_22_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_327 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_22_359 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_22_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_22_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_22_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_22_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_160 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_23_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_324 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_328 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_23_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_23_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_23_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_23_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_23_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_149 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_156 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_24_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_24_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_24_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_24_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_4 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_24_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_24_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_24_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_25_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_25_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_25_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_25_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_25_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_25_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_215 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_291 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_26_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_26_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_26_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_26_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_26_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_26_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_27_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_27_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_27_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_27_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_27_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_27_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_233 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_249 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_28_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_28_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_28_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_28_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_28_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_28_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_112 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_135 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_29_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_306 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_29_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_29_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_29_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_29_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_29_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_29_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_219 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_2_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_2_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_2_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_2_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_2_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_2_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_2_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_113 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_364 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_30_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_30_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_30_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_30_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_30_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_30_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_257 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_31_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_31_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_31_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_31_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_31_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_31_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_120 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_124 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_217 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_223 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_287 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_375 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_32_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_32_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_32_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_32_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_32_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_32_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_147 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_33_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_262 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_289 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_335 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_343 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_347 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_33_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_33_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_33_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_33_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_33_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_33_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_222 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_238 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_299 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_331 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_363 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_383 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_34_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_34_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_34_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_34_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_34_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_34_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_105 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_325 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_35_329 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_35_379 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_35_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_35_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_35_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_35_99 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_123 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_36_225 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_229 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_36_236 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_36_321 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_36_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_36_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_36_86 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_36_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_154 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_37_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_315 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_319 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_37_35 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_37_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_37_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_37_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_37_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_37_92 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_293 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_295 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_356 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_38_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_380 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_38_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_38_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_38_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_38_82 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_38_98 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_152 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_16 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_176 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_26 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_261 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_265 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_273 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_277 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_298 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_310 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_39_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_39_342 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_39_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_39_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_39_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_39_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_39_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_3_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_3_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_3_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_3_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_3_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_3_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_3_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_263 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_290 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_294 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_296 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_303 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_362 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_366 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_40_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_40_43 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_56 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_64 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_40_77 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_40_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_40_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_41_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_41_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_41_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_41_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_78 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_80 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_41_83 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_41_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_41_93 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_116 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_129 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_42_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_358 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_374 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_382 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_42_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_42_47 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_42_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_59 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_42_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_42_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_108 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_169 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_173 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_248 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_252 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_43_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_43_305 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_43_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_43_48 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_43_52 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_43_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_43_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_243 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_253 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_285 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_309 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_313 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_349 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_353 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_357 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_44_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_373 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_44_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_44_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_44_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_44_89 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_44_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_110 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_45_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_45_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_254 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_256 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_286 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_45_316 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_45_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_45_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_45_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_45_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_140 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_148 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_307 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_46_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_337 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_345 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_46_377 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_46_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_46_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_46_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_46_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_100 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_114 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_134 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_138 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_47_175 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_242 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_246 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_250 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_266 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_47_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_47_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_47_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_47_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_47_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_47_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_48_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_143 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_161 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_198 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_202 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_218 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_226 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_230 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_48_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_403 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_41 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_411 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_48_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_48_65 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_48_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_48_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_48_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_179 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_18 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_183 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_190 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_194 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_49_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_234 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_49_268 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_49_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_49_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_49_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_49_74 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_49_96 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_4_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_4_237 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_4_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_4_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_4_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_4_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_111 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_186 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_195 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_207 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_211 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_227 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_235 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_239 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_50_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_50_333 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_341 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_365 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_50_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_50_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_393 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_55 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_50_62 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_50_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_121 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_157 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_241 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_245 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_260 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_272 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_28 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_288 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_32 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_51_320 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_336 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_344 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_348 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_51_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_40 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_46 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_57 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_51_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_51_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_51_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_51_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_102 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_117 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_166 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_193 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_231 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_297 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_301 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_308 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_312 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_33 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_39 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_413 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_417 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_73 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_52_81 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_52_85 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_52_87 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_52_94 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_53_146 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_197 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_205 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_214 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_221 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_259 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_274 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_53_404 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_67 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_69 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_53_76 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_84 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_53_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_53_90 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_53_97 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_104 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_106 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_115 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_127 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_131 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_144 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_151 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_167 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_178 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_187 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_199 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_203 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_206 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_210 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_267 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_300 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_304 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_334 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_338 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_36 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_368 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_372 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_402 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_406 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_410 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_45 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_49 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_51 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_54 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_54_70 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_79 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_54_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_54_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_5_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_136 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_5_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_276 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_5_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_5_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_5_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_5_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_5_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_101 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_155 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_163 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_165 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_172 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_174 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_6_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_189 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_6_220 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_6_224 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_247 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_311 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_6_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_6_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_6_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_6_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_12 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_128 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_132 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_150 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_180 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_184 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_188 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_204 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_216 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_228 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_232 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_264 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_7_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_7_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_384 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_400 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_7_408 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_44 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_7_60 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_68 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_7_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_8 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_7_88 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_91 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_7_95 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_103 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_107 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_118 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_122 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_126 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_130 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_171 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_177 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_181 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_192 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_196 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_2 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_200 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_208 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_22 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_240 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_244 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_278 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_30 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_314 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_8_317 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_34 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_37 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_8_381 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_8_387 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_419 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_8_53 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_8_6 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_8_61 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_8_63 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_32 FILLER_0_9_10 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_119 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_133 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_137 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_139 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_142 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_158 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_164 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_185 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_201 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_209 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_212 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_251 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_255 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_271 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_1 FILLER_0_9_279 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_282 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_346 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_64 FILLER_0_9_352 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_416 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_42 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_8 FILLER_0_9_58 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_4 FILLER_0_9_66 ();
 gf180mcu_fd_sc_mcu7t5v0__fillcap_16 FILLER_0_9_72 ();
 gf180mcu_fd_sc_mcu7t5v0__fill_2 FILLER_0_9_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Left_55 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_0_Right_0 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Left_65 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_10_Right_10 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Left_66 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_11_Right_11 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Left_67 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_12_Right_12 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Left_68 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_13_Right_13 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Left_69 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_14_Right_14 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Left_70 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_15_Right_15 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Left_71 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_16_Right_16 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Left_72 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_17_Right_17 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Left_73 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_18_Right_18 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Left_74 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_19_Right_19 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Left_56 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_1_Right_1 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Left_75 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_20_Right_20 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Left_76 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_21_Right_21 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Left_77 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_22_Right_22 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Left_78 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_23_Right_23 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Left_79 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_24_Right_24 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Left_80 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_25_Right_25 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Left_81 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_26_Right_26 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Left_82 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_27_Right_27 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Left_83 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_28_Right_28 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Left_84 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_29_Right_29 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Left_57 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_2_Right_2 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Left_85 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_30_Right_30 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Left_86 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_31_Right_31 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Left_87 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_32_Right_32 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Left_88 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_33_Right_33 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Left_89 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_34_Right_34 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Left_90 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_35_Right_35 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Left_91 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_36_Right_36 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Left_92 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_37_Right_37 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Left_93 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_38_Right_38 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Left_94 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_39_Right_39 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Left_58 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_3_Right_3 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Left_95 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_40_Right_40 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Left_96 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_41_Right_41 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Left_97 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_42_Right_42 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Left_98 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_43_Right_43 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Left_99 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_44_Right_44 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Left_100 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_45_Right_45 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Left_101 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_46_Right_46 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Left_102 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_47_Right_47 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Left_103 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_48_Right_48 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Left_104 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_49_Right_49 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Left_59 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_4_Right_4 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Left_105 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_50_Right_50 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Left_106 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_51_Right_51 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Left_107 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_52_Right_52 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Left_108 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_53_Right_53 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Left_109 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_54_Right_54 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Left_60 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_5_Right_5 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Left_61 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_6_Right_6 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Left_62 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_7_Right_7 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Left_63 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_8_Right_8 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Left_64 ();
 gf180mcu_fd_sc_mcu7t5v0__endcap PHY_EDGE_ROW_9_Right_9 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_110 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_111 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_112 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_113 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_114 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_115 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_116 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_117 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_118 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_119 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_120 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_0_121 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_171 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_172 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_173 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_174 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_175 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_10_176 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_177 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_178 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_179 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_180 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_11_181 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_182 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_183 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_184 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_185 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_186 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_12_187 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_188 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_189 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_190 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_191 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_13_192 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_193 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_194 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_195 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_196 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_197 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_14_198 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_199 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_200 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_201 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_202 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_15_203 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_204 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_205 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_206 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_207 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_208 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_16_209 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_210 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_211 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_212 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_213 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_17_214 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_215 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_216 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_217 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_218 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_219 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_18_220 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_221 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_222 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_223 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_224 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_19_225 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_122 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_123 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_124 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_125 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_1_126 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_226 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_227 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_228 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_229 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_230 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_20_231 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_232 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_233 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_234 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_235 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_21_236 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_237 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_238 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_239 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_240 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_241 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_22_242 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_243 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_244 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_245 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_246 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_23_247 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_248 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_249 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_250 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_251 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_252 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_24_253 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_254 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_255 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_256 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_257 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_25_258 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_259 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_260 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_261 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_262 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_263 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_26_264 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_265 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_266 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_267 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_268 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_27_269 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_270 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_271 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_272 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_273 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_274 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_28_275 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_276 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_277 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_278 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_279 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_29_280 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_127 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_128 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_129 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_130 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_131 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_2_132 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_281 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_282 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_283 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_284 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_285 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_30_286 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_287 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_288 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_289 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_290 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_31_291 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_292 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_293 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_294 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_295 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_296 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_32_297 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_298 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_299 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_300 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_301 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_33_302 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_303 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_304 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_305 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_306 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_307 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_34_308 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_309 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_310 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_311 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_312 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_35_313 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_314 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_315 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_316 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_317 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_318 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_36_319 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_320 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_321 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_322 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_323 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_37_324 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_325 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_326 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_327 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_328 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_329 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_38_330 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_331 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_332 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_333 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_334 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_39_335 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_133 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_134 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_135 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_136 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_3_137 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_336 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_337 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_338 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_339 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_340 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_40_341 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_342 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_343 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_344 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_345 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_41_346 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_347 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_348 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_349 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_350 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_351 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_42_352 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_353 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_354 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_355 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_356 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_43_357 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_358 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_359 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_360 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_361 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_362 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_44_363 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_364 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_365 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_366 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_367 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_45_368 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_369 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_370 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_371 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_372 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_373 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_46_374 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_375 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_376 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_377 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_378 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_47_379 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_380 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_381 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_382 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_383 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_384 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_48_385 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_386 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_387 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_388 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_389 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_49_390 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_138 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_139 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_140 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_141 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_142 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_4_143 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_391 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_392 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_393 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_394 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_395 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_50_396 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_397 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_398 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_399 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_400 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_51_401 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_402 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_403 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_404 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_405 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_406 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_52_407 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_408 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_409 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_410 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_411 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_53_412 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_413 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_414 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_415 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_416 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_417 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_418 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_419 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_420 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_421 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_422 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_423 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_54_424 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_144 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_145 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_146 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_147 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_5_148 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_149 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_150 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_151 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_152 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_153 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_6_154 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_155 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_156 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_157 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_158 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_7_159 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_160 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_161 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_162 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_163 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_164 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_8_165 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_166 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_167 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_168 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_169 ();
 gf180mcu_fd_sc_mcu7t5v0__filltie TAP_TAPCELL_ROW_9_170 ();
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _400_ (.I(\SPA[0] ),
    .ZN(_070_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _401_ (.A1(_070_),
    .A2(\PORTA[0] ),
    .Z(_071_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _402_ (.I(_071_),
    .Z(net67));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _403_ (.I0(\PORTA[1] ),
    .I1(net5),
    .S(\SPA[1] ),
    .Z(_072_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _404_ (.I(_072_),
    .Z(net74));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _405_ (.I(\SPA[2] ),
    .ZN(_073_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _406_ (.A1(_073_),
    .A2(\PORTA[2] ),
    .Z(_074_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _407_ (.I(_074_),
    .Z(net75));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _408_ (.I0(\PORTA[3] ),
    .I1(net40),
    .S(\SPA[3] ),
    .Z(_075_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _409_ (.I(_075_),
    .Z(net76));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _410_ (.I0(\PORTA[4] ),
    .I1(net41),
    .S(\SPA[4] ),
    .Z(_076_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _411_ (.I(_076_),
    .Z(net77));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _412_ (.I0(\PORTA[5] ),
    .I1(net36),
    .S(\SPA[5] ),
    .Z(_077_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _413_ (.I(_077_),
    .Z(net78));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _414_ (.I0(\PORTA[6] ),
    .I1(net37),
    .S(\SPA[6] ),
    .Z(_078_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _415_ (.I(_078_),
    .Z(net79));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _416_ (.I(\SPA[7] ),
    .ZN(_079_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _417_ (.A1(_079_),
    .A2(\PORTA[7] ),
    .Z(_080_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _418_ (.I(_080_),
    .Z(net80));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _419_ (.A1(\SPA[1] ),
    .A2(\DDRA[1] ),
    .ZN(net58));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _420_ (.A1(\SPA[3] ),
    .A2(\DDRA[3] ),
    .ZN(net60));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _421_ (.A1(\SPA[4] ),
    .A2(\DDRA[4] ),
    .ZN(net61));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _422_ (.A1(\SPA[5] ),
    .A2(\DDRA[5] ),
    .ZN(net62));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _423_ (.A1(\SPA[6] ),
    .A2(\DDRA[6] ),
    .ZN(net63));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _424_ (.I(net28),
    .ZN(_081_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _425_ (.A1(\SPA[2] ),
    .A2(_081_),
    .ZN(net42));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _426_ (.I(\SPB[0] ),
    .ZN(_082_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _427_ (.A1(_082_),
    .A2(\PORTB[0] ),
    .Z(_083_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _428_ (.I(_083_),
    .Z(net81));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _429_ (.I0(\PORTB[1] ),
    .I1(net38),
    .S(\SPB[1] ),
    .Z(_084_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _430_ (.I(_084_),
    .Z(net82));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _431_ (.I(\SPB[2] ),
    .Z(_085_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _432_ (.I(\PORTB[2] ),
    .ZN(_086_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _433_ (.A1(_085_),
    .A2(_086_),
    .ZN(net68));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _434_ (.I(\SPB[3] ),
    .ZN(_087_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _435_ (.A1(_087_),
    .A2(\PORTB[3] ),
    .Z(_088_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _436_ (.I(_088_),
    .Z(net69));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _437_ (.I0(\PORTB[4] ),
    .I1(net3),
    .S(\SPB[4] ),
    .Z(_089_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _438_ (.I(_089_),
    .Z(net70));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _439_ (.I0(\PORTB[5] ),
    .I1(net2),
    .S(\SPB[5] ),
    .Z(_090_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _440_ (.I(_090_),
    .Z(net71));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _441_ (.I0(\PORTB[6] ),
    .I1(net4),
    .S(\SPB[6] ),
    .Z(_091_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _442_ (.I(_091_),
    .Z(net72));
 gf180mcu_fd_sc_mcu7t5v0__mux2_2 _443_ (.I0(\PORTB[7] ),
    .I1(net1),
    .S(\SPB[7] ),
    .Z(_092_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _444_ (.I(_092_),
    .Z(net73));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _445_ (.A1(\SPB[1] ),
    .A2(\DDRB[1] ),
    .ZN(net66));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _446_ (.A1(\SPB[4] ),
    .A2(\DDRB[4] ),
    .ZN(net54));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _447_ (.A1(\SPB[5] ),
    .A2(\DDRB[5] ),
    .ZN(net55));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _448_ (.A1(\SPB[6] ),
    .A2(\DDRB[6] ),
    .ZN(net56));
 gf180mcu_fd_sc_mcu7t5v0__nor2_2 _449_ (.A1(\SPB[7] ),
    .A2(\DDRB[7] ),
    .ZN(net57));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _450_ (.A1(_070_),
    .A2(\DDRA[0] ),
    .ZN(net51));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _451_ (.A1(_073_),
    .A2(\DDRA[2] ),
    .ZN(net59));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _452_ (.A1(_079_),
    .A2(\DDRA[7] ),
    .ZN(net64));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _453_ (.A1(_082_),
    .A2(\DDRB[0] ),
    .ZN(net65));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _454_ (.I(\DDRB[2] ),
    .ZN(_093_));
 gf180mcu_fd_sc_mcu7t5v0__or2_1 _455_ (.A1(_085_),
    .A2(_093_),
    .Z(_094_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _456_ (.I(_094_),
    .Z(net52));
 gf180mcu_fd_sc_mcu7t5v0__nand2_2 _457_ (.A1(_087_),
    .A2(\DDRB[3] ),
    .ZN(net53));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _458_ (.A1(_085_),
    .A2(net21),
    .Z(_095_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _459_ (.I(_095_),
    .Z(net94));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _460_ (.A1(\SPB[3] ),
    .A2(net22),
    .Z(_096_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _461_ (.I(_096_),
    .Z(net95));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _462_ (.I(net39),
    .Z(_097_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _463_ (.I(_097_),
    .Z(_098_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _464_ (.I(_098_),
    .Z(_099_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _465_ (.A1(\SPA[7] ),
    .A2(net33),
    .ZN(_100_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _466_ (.A1(_099_),
    .A2(_100_),
    .ZN(_000_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _467_ (.I(net10),
    .Z(_101_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _468_ (.I(_101_),
    .ZN(_102_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _469_ (.I(_102_),
    .Z(_103_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _470_ (.I(_103_),
    .Z(_104_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _471_ (.I(net43),
    .ZN(_105_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _472_ (.I(net9),
    .Z(_106_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _473_ (.I(net6),
    .Z(_107_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _474_ (.I(net7),
    .Z(_108_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_1 _475_ (.A1(_107_),
    .A2(_108_),
    .A3(net8),
    .ZN(_109_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _476_ (.A1(_106_),
    .A2(_109_),
    .Z(_110_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _477_ (.I(_110_),
    .Z(_111_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _478_ (.I(net6),
    .ZN(_112_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 _479_ (.I(_112_),
    .Z(_113_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_3 _480_ (.I(net7),
    .ZN(_114_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _481_ (.I(_114_),
    .Z(_115_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_2 _482_ (.I(net8),
    .ZN(_116_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _483_ (.I(_116_),
    .Z(_117_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _484_ (.I(net9),
    .Z(_118_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _485_ (.A1(_113_),
    .A2(_115_),
    .A3(_117_),
    .A4(_118_),
    .ZN(_119_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _486_ (.I(_119_),
    .Z(_120_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _487_ (.I(_108_),
    .Z(_121_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _488_ (.A1(_113_),
    .A2(_121_),
    .A3(_117_),
    .A4(_118_),
    .ZN(_122_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _489_ (.I(_122_),
    .Z(_123_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _490_ (.A1(\SPB[0] ),
    .A2(_111_),
    .B1(_120_),
    .B2(net83),
    .C1(_123_),
    .C2(net20),
    .ZN(_124_));
 gf180mcu_fd_sc_mcu7t5v0__or2_2 _491_ (.A1(net8),
    .A2(_106_),
    .Z(_125_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _492_ (.A1(_113_),
    .A2(_121_),
    .A3(_125_),
    .ZN(_126_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _493_ (.A1(_112_),
    .A2(_114_),
    .A3(_125_),
    .ZN(_127_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _494_ (.I(_127_),
    .Z(_128_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _495_ (.A1(\DDRB[0] ),
    .A2(_126_),
    .B1(_128_),
    .B2(\PORTB[0] ),
    .ZN(_129_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _496_ (.I(net8),
    .Z(_130_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _497_ (.I(net9),
    .ZN(_131_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _498_ (.A1(_112_),
    .A2(_108_),
    .A3(_130_),
    .A4(_131_),
    .ZN(_132_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _499_ (.I(_132_),
    .Z(_133_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _500_ (.I(_107_),
    .Z(_134_));
 gf180mcu_fd_sc_mcu7t5v0__nor3_4 _501_ (.A1(_134_),
    .A2(_114_),
    .A3(_125_),
    .ZN(_135_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _502_ (.I(_135_),
    .Z(_136_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _503_ (.A1(_107_),
    .A2(_108_),
    .A3(_116_),
    .A4(_106_),
    .ZN(_137_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _504_ (.I(_137_),
    .Z(_138_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _505_ (.A1(net86),
    .A2(_133_),
    .B1(_136_),
    .B2(\PORTA[0] ),
    .C1(\SPA[0] ),
    .C2(_138_),
    .ZN(_139_));
 gf180mcu_fd_sc_mcu7t5v0__nor4_4 _506_ (.A1(_107_),
    .A2(_114_),
    .A3(_116_),
    .A4(_106_),
    .ZN(_140_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _507_ (.I(_131_),
    .Z(_141_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _508_ (.A1(_141_),
    .A2(_109_),
    .Z(_142_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _509_ (.I(_142_),
    .Z(_143_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _510_ (.I(_102_),
    .Z(_144_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _511_ (.A1(net34),
    .A2(_140_),
    .B1(_143_),
    .B2(\DDRA[0] ),
    .C(_144_),
    .ZN(_145_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _512_ (.A1(_129_),
    .A2(_139_),
    .A3(_145_),
    .Z(_146_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _513_ (.I(_097_),
    .Z(_147_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _514_ (.A1(_104_),
    .A2(_105_),
    .B1(_124_),
    .B2(_146_),
    .C(_147_),
    .ZN(_001_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _515_ (.I(net44),
    .ZN(_148_));
 gf180mcu_fd_sc_mcu7t5v0__oai21_2 _516_ (.A1(_121_),
    .A2(_130_),
    .B(_118_),
    .ZN(_149_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _517_ (.A1(\DDRB[1] ),
    .A2(_126_),
    .B1(_143_),
    .B2(\DDRA[1] ),
    .ZN(_150_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _518_ (.A1(_149_),
    .A2(_150_),
    .Z(_151_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _519_ (.A1(net35),
    .A2(_140_),
    .B1(_136_),
    .B2(\PORTA[1] ),
    .C1(\SPA[1] ),
    .C2(_138_),
    .ZN(_152_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _520_ (.A1(net87),
    .A2(_133_),
    .B1(_122_),
    .B2(net27),
    .C(_144_),
    .ZN(_153_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _521_ (.I(_110_),
    .Z(_154_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _522_ (.I(_127_),
    .Z(_155_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _523_ (.A1(\SPB[1] ),
    .A2(_154_),
    .B1(_155_),
    .B2(\PORTB[1] ),
    .ZN(_156_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _524_ (.A1(_152_),
    .A2(_153_),
    .A3(_156_),
    .Z(_157_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _525_ (.A1(_104_),
    .A2(_148_),
    .B1(_151_),
    .B2(_157_),
    .C(_147_),
    .ZN(_002_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _526_ (.I(net45),
    .ZN(_158_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_4 _527_ (.A1(_134_),
    .A2(_115_),
    .A3(_117_),
    .A4(_141_),
    .ZN(_159_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _528_ (.A1(_134_),
    .A2(_115_),
    .A3(_130_),
    .A4(_141_),
    .ZN(_160_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _529_ (.A1(_093_),
    .A2(_159_),
    .B1(_160_),
    .B2(_081_),
    .ZN(_161_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _530_ (.A1(\SPB[2] ),
    .A2(_111_),
    .B1(_155_),
    .B2(\PORTB[2] ),
    .C(_161_),
    .ZN(_162_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _531_ (.I(_140_),
    .Z(_163_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _532_ (.I(_132_),
    .Z(_164_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _533_ (.I(_137_),
    .Z(_165_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _534_ (.A1(net21),
    .A2(_163_),
    .B1(_164_),
    .B2(net88),
    .C1(\SPA[2] ),
    .C2(_165_),
    .ZN(_166_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _535_ (.I(_135_),
    .Z(_167_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _536_ (.A1(\PORTA[2] ),
    .A2(_167_),
    .B1(_143_),
    .B2(\DDRA[2] ),
    .C(_103_),
    .ZN(_168_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _537_ (.A1(_166_),
    .A2(_168_),
    .Z(_169_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _538_ (.I(_097_),
    .Z(_170_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _539_ (.A1(_104_),
    .A2(_158_),
    .B1(_162_),
    .B2(_169_),
    .C(_170_),
    .ZN(_003_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _540_ (.I(_103_),
    .Z(_171_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _541_ (.I(net46),
    .ZN(_172_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _542_ (.I(_126_),
    .Z(_173_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _543_ (.I(_142_),
    .Z(_174_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _544_ (.A1(\SPB[3] ),
    .A2(_111_),
    .B1(_173_),
    .B2(\DDRB[3] ),
    .C1(_174_),
    .C2(\DDRA[3] ),
    .ZN(_175_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _545_ (.A1(net22),
    .A2(_140_),
    .B1(_135_),
    .B2(\PORTA[3] ),
    .C1(\SPA[3] ),
    .C2(_138_),
    .ZN(_176_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _546_ (.A1(\PORTB[3] ),
    .A2(_128_),
    .B1(_122_),
    .B2(net29),
    .ZN(_177_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _547_ (.A1(net89),
    .A2(_164_),
    .B(_103_),
    .ZN(_178_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _548_ (.A1(_149_),
    .A2(_176_),
    .A3(_177_),
    .A4(_178_),
    .Z(_179_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _549_ (.A1(_171_),
    .A2(_172_),
    .B1(_175_),
    .B2(_179_),
    .C(_170_),
    .ZN(_004_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _550_ (.I(net47),
    .ZN(_180_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _551_ (.I(\DDRB[4] ),
    .ZN(_181_));
 gf180mcu_fd_sc_mcu7t5v0__inv_1 _552_ (.I(net30),
    .ZN(_182_));
 gf180mcu_fd_sc_mcu7t5v0__oai22_1 _553_ (.A1(_181_),
    .A2(_159_),
    .B1(_160_),
    .B2(_182_),
    .ZN(_183_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _554_ (.A1(\PORTB[4] ),
    .A2(_155_),
    .B1(_174_),
    .B2(\DDRA[4] ),
    .C(_183_),
    .ZN(_184_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_1 _555_ (.A1(net90),
    .A2(_133_),
    .B1(_167_),
    .B2(\PORTA[4] ),
    .C1(\SPA[4] ),
    .C2(_165_),
    .ZN(_185_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _556_ (.A1(\SPB[4] ),
    .A2(_111_),
    .B1(_163_),
    .B2(net23),
    .C(_144_),
    .ZN(_186_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _557_ (.A1(_185_),
    .A2(_186_),
    .Z(_187_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _558_ (.A1(_171_),
    .A2(_180_),
    .B1(_184_),
    .B2(_187_),
    .C(_170_),
    .ZN(_005_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _559_ (.I(net48),
    .ZN(_188_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _560_ (.A1(\DDRB[5] ),
    .A2(_173_),
    .B1(_174_),
    .B2(\DDRA[5] ),
    .C1(_155_),
    .C2(\PORTB[5] ),
    .ZN(_189_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _561_ (.A1(_101_),
    .A2(_149_),
    .Z(_190_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _562_ (.A1(\PORTA[5] ),
    .A2(_167_),
    .B1(_165_),
    .B2(\SPA[5] ),
    .ZN(_191_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _563_ (.A1(net24),
    .A2(_163_),
    .B1(_164_),
    .B2(net91),
    .ZN(_192_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _564_ (.A1(\SPB[5] ),
    .A2(_154_),
    .B1(_123_),
    .B2(net31),
    .ZN(_193_));
 gf180mcu_fd_sc_mcu7t5v0__and4_1 _565_ (.A1(_190_),
    .A2(_191_),
    .A3(_192_),
    .A4(_193_),
    .Z(_194_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _566_ (.A1(_171_),
    .A2(_188_),
    .B1(_189_),
    .B2(_194_),
    .C(_170_),
    .ZN(_006_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _567_ (.I(net49),
    .ZN(_195_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _568_ (.A1(\DDRB[6] ),
    .A2(_173_),
    .B1(_174_),
    .B2(\DDRA[6] ),
    .C1(_123_),
    .C2(net32),
    .ZN(_196_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _569_ (.A1(net92),
    .A2(_133_),
    .B1(_136_),
    .B2(\PORTA[6] ),
    .C1(\SPA[6] ),
    .C2(_138_),
    .ZN(_197_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _570_ (.A1(\SPB[6] ),
    .A2(_154_),
    .B1(_163_),
    .B2(net25),
    .C(_144_),
    .ZN(_198_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _571_ (.A1(\PORTB[6] ),
    .A2(_128_),
    .B1(_119_),
    .B2(net84),
    .ZN(_199_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _572_ (.A1(_197_),
    .A2(_198_),
    .A3(_199_),
    .Z(_200_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _573_ (.A1(_171_),
    .A2(_195_),
    .B1(_196_),
    .B2(_200_),
    .C(_098_),
    .ZN(_007_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _574_ (.I(net50),
    .ZN(_201_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _575_ (.I(net26),
    .ZN(_202_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_2 _576_ (.A1(_113_),
    .A2(_121_),
    .A3(_130_),
    .A4(_141_),
    .ZN(_203_));
 gf180mcu_fd_sc_mcu7t5v0__oai211_2 _577_ (.A1(_202_),
    .A2(_203_),
    .B(_149_),
    .C(_101_),
    .ZN(_204_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_2 _578_ (.A1(\DDRB[7] ),
    .A2(_173_),
    .B1(_123_),
    .B2(net33),
    .C(_204_),
    .ZN(_205_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _579_ (.A1(net93),
    .A2(_164_),
    .B1(_165_),
    .B2(\SPA[7] ),
    .ZN(_206_));
 gf180mcu_fd_sc_mcu7t5v0__aoi22_1 _580_ (.A1(net85),
    .A2(_119_),
    .B1(_143_),
    .B2(\DDRA[7] ),
    .ZN(_207_));
 gf180mcu_fd_sc_mcu7t5v0__aoi222_2 _581_ (.A1(\SPB[7] ),
    .A2(_154_),
    .B1(_128_),
    .B2(\PORTB[7] ),
    .C1(_167_),
    .C2(\PORTA[7] ),
    .ZN(_208_));
 gf180mcu_fd_sc_mcu7t5v0__and3_1 _582_ (.A1(_206_),
    .A2(_207_),
    .A3(_208_),
    .Z(_209_));
 gf180mcu_fd_sc_mcu7t5v0__aoi221_1 _583_ (.A1(_201_),
    .A2(_104_),
    .B1(_205_),
    .B2(_209_),
    .C(_098_),
    .ZN(_008_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _584_ (.I(net12),
    .Z(_210_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _585_ (.A1(net10),
    .A2(net11),
    .Z(_211_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _586_ (.I(_211_),
    .Z(_212_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _587_ (.I(_212_),
    .Z(_213_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _588_ (.A1(_210_),
    .A2(_120_),
    .A3(_213_),
    .ZN(_214_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _589_ (.A1(\SPA[0] ),
    .A2(net20),
    .ZN(_215_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _590_ (.A1(last_irq0_trigger),
    .A2(_215_),
    .ZN(_216_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _591_ (.A1(net83),
    .A2(_214_),
    .B(_216_),
    .ZN(_217_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _592_ (.A1(_099_),
    .A2(_217_),
    .ZN(_009_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _593_ (.I(net18),
    .Z(_218_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _594_ (.A1(_218_),
    .A2(_120_),
    .A3(_213_),
    .ZN(_219_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _595_ (.A1(\SPB[0] ),
    .A2(net34),
    .ZN(_220_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _596_ (.A1(last_irg6_trigger),
    .A2(_220_),
    .ZN(_221_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _597_ (.A1(net84),
    .A2(_219_),
    .B(_221_),
    .ZN(_222_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _598_ (.A1(_099_),
    .A2(_222_),
    .ZN(_010_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _599_ (.I(net19),
    .Z(_223_));
 gf180mcu_fd_sc_mcu7t5v0__nand3_1 _600_ (.A1(_223_),
    .A2(_120_),
    .A3(_213_),
    .ZN(_224_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _601_ (.A1(last_irq7_trigger),
    .A2(_100_),
    .ZN(_225_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _602_ (.A1(net85),
    .A2(_224_),
    .B(_225_),
    .ZN(_226_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _603_ (.A1(_099_),
    .A2(_226_),
    .ZN(_011_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _604_ (.I(net12),
    .Z(_227_));
 gf180mcu_fd_sc_mcu7t5v0__nand4_1 _605_ (.A1(_134_),
    .A2(_115_),
    .A3(_117_),
    .A4(_118_),
    .ZN(_228_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _606_ (.A1(_101_),
    .A2(net11),
    .ZN(_229_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _607_ (.A1(_228_),
    .A2(_229_),
    .ZN(_230_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _608_ (.I(_230_),
    .Z(_231_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _609_ (.A1(_227_),
    .A2(_231_),
    .ZN(_232_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _610_ (.I(_211_),
    .Z(_233_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _611_ (.A1(_132_),
    .A2(_233_),
    .ZN(_234_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _612_ (.I(_234_),
    .Z(_235_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _613_ (.I(_235_),
    .Z(_236_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _614_ (.A1(net86),
    .A2(_236_),
    .ZN(_237_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _615_ (.I(_098_),
    .Z(_238_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _616_ (.A1(_232_),
    .A2(_237_),
    .B(_238_),
    .ZN(_012_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _617_ (.I(net87),
    .ZN(_239_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _618_ (.A1(net13),
    .A2(_235_),
    .ZN(_240_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _619_ (.I(_097_),
    .Z(_241_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _620_ (.A1(_239_),
    .A2(_236_),
    .B(_240_),
    .C(_241_),
    .ZN(_013_));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 _621_ (.I(net14),
    .Z(_242_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _622_ (.A1(_242_),
    .A2(_231_),
    .ZN(_243_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _623_ (.I(_234_),
    .Z(_244_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _624_ (.A1(net88),
    .A2(_244_),
    .ZN(_245_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _625_ (.A1(_243_),
    .A2(_245_),
    .B(_238_),
    .ZN(_014_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _626_ (.I(net89),
    .ZN(_246_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _627_ (.A1(net15),
    .A2(_235_),
    .ZN(_247_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _628_ (.A1(_246_),
    .A2(_236_),
    .B(_247_),
    .C(_241_),
    .ZN(_015_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _629_ (.I(net16),
    .Z(_248_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _630_ (.A1(_248_),
    .A2(_231_),
    .ZN(_249_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _631_ (.A1(net90),
    .A2(_244_),
    .ZN(_250_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _632_ (.A1(_249_),
    .A2(_250_),
    .B(_238_),
    .ZN(_016_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _633_ (.I(net91),
    .ZN(_251_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _634_ (.A1(net17),
    .A2(_235_),
    .ZN(_252_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _635_ (.I(net39),
    .Z(_253_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _636_ (.I(_253_),
    .Z(_254_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _637_ (.A1(_251_),
    .A2(_236_),
    .B(_252_),
    .C(_254_),
    .ZN(_017_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _638_ (.I(net18),
    .Z(_255_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _639_ (.A1(_255_),
    .A2(_231_),
    .ZN(_256_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _640_ (.A1(net92),
    .A2(_244_),
    .ZN(_257_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _641_ (.A1(_256_),
    .A2(_257_),
    .B(_238_),
    .ZN(_018_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _642_ (.I(net19),
    .Z(_258_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _643_ (.A1(_258_),
    .A2(_230_),
    .ZN(_259_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _644_ (.A1(net93),
    .A2(_244_),
    .ZN(_260_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _645_ (.I(net39),
    .Z(_261_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _646_ (.I(_261_),
    .Z(_262_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _647_ (.A1(_259_),
    .A2(_260_),
    .B(_262_),
    .ZN(_019_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _648_ (.I(_211_),
    .Z(_263_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _649_ (.A1(_142_),
    .A2(_263_),
    .Z(_264_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _650_ (.I(_264_),
    .Z(_265_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _651_ (.A1(_227_),
    .A2(_265_),
    .ZN(_266_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _652_ (.A1(_142_),
    .A2(_213_),
    .ZN(_267_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _653_ (.I(_267_),
    .Z(_268_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _654_ (.A1(\DDRA[0] ),
    .A2(_268_),
    .ZN(_269_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _655_ (.A1(_266_),
    .A2(_269_),
    .B(_262_),
    .ZN(_020_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _656_ (.I(net13),
    .Z(_270_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _657_ (.A1(_270_),
    .A2(_265_),
    .ZN(_271_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _658_ (.A1(\DDRA[1] ),
    .A2(_268_),
    .ZN(_272_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _659_ (.A1(_271_),
    .A2(_272_),
    .B(_262_),
    .ZN(_021_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _660_ (.A1(_242_),
    .A2(_265_),
    .ZN(_273_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _661_ (.A1(\DDRA[2] ),
    .A2(_268_),
    .ZN(_274_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _662_ (.A1(_273_),
    .A2(_274_),
    .B(_262_),
    .ZN(_022_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _663_ (.I(net15),
    .Z(_275_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _664_ (.A1(_275_),
    .A2(_265_),
    .ZN(_276_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _665_ (.A1(\DDRA[3] ),
    .A2(_268_),
    .ZN(_277_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _666_ (.I(_261_),
    .Z(_278_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _667_ (.A1(_276_),
    .A2(_277_),
    .B(_278_),
    .ZN(_023_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _668_ (.I(_264_),
    .Z(_279_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _669_ (.A1(_248_),
    .A2(_279_),
    .ZN(_280_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _670_ (.I(_267_),
    .Z(_281_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _671_ (.A1(\DDRA[4] ),
    .A2(_281_),
    .ZN(_282_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _672_ (.A1(_280_),
    .A2(_282_),
    .B(_278_),
    .ZN(_024_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _673_ (.I(net17),
    .Z(_283_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _674_ (.A1(_283_),
    .A2(_279_),
    .ZN(_284_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _675_ (.A1(\DDRA[5] ),
    .A2(_281_),
    .ZN(_285_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _676_ (.A1(_284_),
    .A2(_285_),
    .B(_278_),
    .ZN(_025_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _677_ (.A1(_255_),
    .A2(_279_),
    .ZN(_286_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _678_ (.A1(\DDRA[6] ),
    .A2(_281_),
    .ZN(_287_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _679_ (.A1(_286_),
    .A2(_287_),
    .B(_278_),
    .ZN(_026_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _680_ (.A1(_258_),
    .A2(_279_),
    .ZN(_288_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _681_ (.A1(\DDRA[7] ),
    .A2(_281_),
    .ZN(_289_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _682_ (.I(_261_),
    .Z(_290_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _683_ (.A1(_288_),
    .A2(_289_),
    .B(_290_),
    .ZN(_027_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _684_ (.A1(_159_),
    .A2(_229_),
    .ZN(_291_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _685_ (.I(_291_),
    .Z(_292_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _686_ (.A1(_227_),
    .A2(_292_),
    .ZN(_293_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _687_ (.A1(_126_),
    .A2(_212_),
    .ZN(_294_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _688_ (.I(_294_),
    .Z(_295_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _689_ (.I(_295_),
    .Z(_296_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _690_ (.A1(\DDRB[0] ),
    .A2(_296_),
    .ZN(_297_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _691_ (.A1(_293_),
    .A2(_297_),
    .B(_290_),
    .ZN(_028_));
 gf180mcu_fd_sc_mcu7t5v0__clkinv_1 _692_ (.I(\DDRB[1] ),
    .ZN(_298_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _693_ (.A1(net13),
    .A2(_295_),
    .ZN(_299_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _694_ (.A1(_298_),
    .A2(_296_),
    .B(_299_),
    .C(_254_),
    .ZN(_029_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _695_ (.A1(net14),
    .A2(_295_),
    .ZN(_300_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _696_ (.A1(_093_),
    .A2(_296_),
    .B(_300_),
    .C(_254_),
    .ZN(_030_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _697_ (.A1(_275_),
    .A2(_292_),
    .ZN(_301_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _698_ (.I(_294_),
    .Z(_302_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _699_ (.A1(\DDRB[3] ),
    .A2(_302_),
    .ZN(_303_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _700_ (.A1(_301_),
    .A2(_303_),
    .B(_290_),
    .ZN(_031_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _701_ (.A1(net16),
    .A2(_295_),
    .ZN(_304_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _702_ (.A1(_181_),
    .A2(_296_),
    .B(_304_),
    .C(_254_),
    .ZN(_032_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _703_ (.A1(_283_),
    .A2(_292_),
    .ZN(_305_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _704_ (.A1(\DDRB[5] ),
    .A2(_302_),
    .ZN(_306_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _705_ (.A1(_305_),
    .A2(_306_),
    .B(_290_),
    .ZN(_033_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _706_ (.A1(_255_),
    .A2(_292_),
    .ZN(_307_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _707_ (.A1(\DDRB[6] ),
    .A2(_302_),
    .ZN(_308_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 _708_ (.I(_261_),
    .Z(_309_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _709_ (.A1(_307_),
    .A2(_308_),
    .B(_309_),
    .ZN(_034_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _710_ (.A1(_258_),
    .A2(_291_),
    .ZN(_310_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _711_ (.A1(\DDRB[7] ),
    .A2(_302_),
    .ZN(_311_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _712_ (.A1(_310_),
    .A2(_311_),
    .B(_309_),
    .ZN(_035_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _713_ (.A1(_135_),
    .A2(_263_),
    .Z(_312_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _714_ (.I(_312_),
    .Z(_313_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _715_ (.A1(_227_),
    .A2(_313_),
    .ZN(_314_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _716_ (.A1(_136_),
    .A2(_263_),
    .ZN(_315_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _717_ (.I(_315_),
    .Z(_316_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _718_ (.A1(\PORTA[0] ),
    .A2(_316_),
    .ZN(_317_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _719_ (.A1(_314_),
    .A2(_317_),
    .B(_309_),
    .ZN(_036_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _720_ (.A1(_270_),
    .A2(_313_),
    .ZN(_318_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _721_ (.A1(\PORTA[1] ),
    .A2(_316_),
    .ZN(_319_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _722_ (.A1(_318_),
    .A2(_319_),
    .B(_309_),
    .ZN(_037_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _723_ (.A1(_242_),
    .A2(_313_),
    .ZN(_320_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _724_ (.A1(\PORTA[2] ),
    .A2(_316_),
    .ZN(_321_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _725_ (.I(net39),
    .Z(_322_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _726_ (.I(_322_),
    .Z(_323_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _727_ (.A1(_320_),
    .A2(_321_),
    .B(_323_),
    .ZN(_038_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _728_ (.A1(_275_),
    .A2(_313_),
    .ZN(_324_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _729_ (.A1(\PORTA[3] ),
    .A2(_316_),
    .ZN(_325_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _730_ (.A1(_324_),
    .A2(_325_),
    .B(_323_),
    .ZN(_039_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _731_ (.I(_312_),
    .Z(_326_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _732_ (.A1(_248_),
    .A2(_326_),
    .ZN(_327_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _733_ (.I(_315_),
    .Z(_328_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _734_ (.A1(\PORTA[4] ),
    .A2(_328_),
    .ZN(_329_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _735_ (.A1(_327_),
    .A2(_329_),
    .B(_323_),
    .ZN(_040_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _736_ (.A1(_283_),
    .A2(_326_),
    .ZN(_330_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _737_ (.A1(\PORTA[5] ),
    .A2(_328_),
    .ZN(_331_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _738_ (.A1(_330_),
    .A2(_331_),
    .B(_323_),
    .ZN(_041_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _739_ (.A1(_255_),
    .A2(_326_),
    .ZN(_332_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _740_ (.A1(\PORTA[6] ),
    .A2(_328_),
    .ZN(_333_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _741_ (.I(_322_),
    .Z(_334_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _742_ (.A1(_332_),
    .A2(_333_),
    .B(_334_),
    .ZN(_042_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _743_ (.A1(_258_),
    .A2(_326_),
    .ZN(_335_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _744_ (.A1(\PORTA[7] ),
    .A2(_328_),
    .ZN(_336_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _745_ (.A1(_335_),
    .A2(_336_),
    .B(_334_),
    .ZN(_043_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _746_ (.A1(_127_),
    .A2(_233_),
    .Z(_337_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _747_ (.I(_337_),
    .Z(_338_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _748_ (.A1(_210_),
    .A2(_338_),
    .ZN(_339_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _749_ (.A1(_127_),
    .A2(_212_),
    .ZN(_340_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _750_ (.I(_340_),
    .Z(_341_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _751_ (.A1(\PORTB[0] ),
    .A2(_341_),
    .ZN(_342_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _752_ (.A1(_339_),
    .A2(_342_),
    .B(_334_),
    .ZN(_044_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _753_ (.A1(_270_),
    .A2(_338_),
    .ZN(_343_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _754_ (.A1(\PORTB[1] ),
    .A2(_341_),
    .ZN(_344_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _755_ (.A1(_343_),
    .A2(_344_),
    .B(_334_),
    .ZN(_045_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _756_ (.A1(net14),
    .A2(_340_),
    .ZN(_345_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _757_ (.I(_253_),
    .Z(_346_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _758_ (.A1(_086_),
    .A2(_341_),
    .B(_345_),
    .C(_346_),
    .ZN(_046_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _759_ (.A1(_275_),
    .A2(_338_),
    .ZN(_347_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _760_ (.A1(\PORTB[3] ),
    .A2(_341_),
    .ZN(_348_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _761_ (.I(_322_),
    .Z(_349_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _762_ (.A1(_347_),
    .A2(_348_),
    .B(_349_),
    .ZN(_047_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _763_ (.A1(_248_),
    .A2(_338_),
    .ZN(_350_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _764_ (.I(_340_),
    .Z(_351_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _765_ (.A1(\PORTB[4] ),
    .A2(_351_),
    .ZN(_352_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _766_ (.A1(_350_),
    .A2(_352_),
    .B(_349_),
    .ZN(_048_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _767_ (.A1(_283_),
    .A2(_337_),
    .ZN(_353_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _768_ (.A1(\PORTB[5] ),
    .A2(_351_),
    .ZN(_354_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _769_ (.A1(_353_),
    .A2(_354_),
    .B(_349_),
    .ZN(_049_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _770_ (.A1(_218_),
    .A2(_337_),
    .ZN(_355_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _771_ (.A1(\PORTB[6] ),
    .A2(_351_),
    .ZN(_356_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _772_ (.A1(_355_),
    .A2(_356_),
    .B(_349_),
    .ZN(_050_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _773_ (.A1(_223_),
    .A2(_337_),
    .ZN(_357_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _774_ (.A1(\PORTB[7] ),
    .A2(_351_),
    .ZN(_358_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _775_ (.I(_322_),
    .Z(_359_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _776_ (.A1(_357_),
    .A2(_358_),
    .B(_359_),
    .ZN(_051_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _777_ (.A1(_137_),
    .A2(_212_),
    .ZN(_360_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _778_ (.I(_360_),
    .Z(_361_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _779_ (.I(_361_),
    .Z(_362_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _780_ (.A1(_210_),
    .A2(_361_),
    .ZN(_363_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _781_ (.A1(_070_),
    .A2(_362_),
    .B(_363_),
    .C(_346_),
    .ZN(_052_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _782_ (.A1(_137_),
    .A2(_233_),
    .Z(_364_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _783_ (.I(_364_),
    .Z(_365_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _784_ (.A1(_270_),
    .A2(_365_),
    .ZN(_366_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _785_ (.A1(\SPA[1] ),
    .A2(_362_),
    .ZN(_367_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _786_ (.A1(_366_),
    .A2(_367_),
    .B(_359_),
    .ZN(_053_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _787_ (.A1(net14),
    .A2(_361_),
    .ZN(_368_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _788_ (.A1(_073_),
    .A2(_362_),
    .B(_368_),
    .C(_346_),
    .ZN(_054_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _789_ (.A1(net15),
    .A2(_365_),
    .ZN(_369_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _790_ (.I(_360_),
    .Z(_370_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _791_ (.A1(\SPA[3] ),
    .A2(_370_),
    .ZN(_371_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _792_ (.A1(_369_),
    .A2(_371_),
    .B(_359_),
    .ZN(_055_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _793_ (.A1(net16),
    .A2(_365_),
    .ZN(_372_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _794_ (.A1(\SPA[4] ),
    .A2(_370_),
    .ZN(_373_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _795_ (.A1(_372_),
    .A2(_373_),
    .B(_359_),
    .ZN(_056_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _796_ (.A1(net17),
    .A2(_365_),
    .ZN(_374_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _797_ (.A1(\SPA[5] ),
    .A2(_370_),
    .ZN(_375_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _798_ (.I(_253_),
    .Z(_376_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _799_ (.A1(_374_),
    .A2(_375_),
    .B(_376_),
    .ZN(_057_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _800_ (.A1(_218_),
    .A2(_364_),
    .ZN(_377_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _801_ (.A1(\SPA[6] ),
    .A2(_370_),
    .ZN(_378_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _802_ (.A1(_377_),
    .A2(_378_),
    .B(_376_),
    .ZN(_058_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _803_ (.A1(_223_),
    .A2(_361_),
    .ZN(_379_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _804_ (.A1(_079_),
    .A2(_362_),
    .B(_379_),
    .C(_346_),
    .ZN(_059_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _805_ (.A1(_110_),
    .A2(_263_),
    .ZN(_380_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _806_ (.I(_380_),
    .Z(_381_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _807_ (.A1(_210_),
    .A2(_380_),
    .ZN(_382_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _808_ (.A1(_082_),
    .A2(_381_),
    .B(_382_),
    .C(_147_),
    .ZN(_060_));
 gf180mcu_fd_sc_mcu7t5v0__and2_1 _809_ (.A1(_110_),
    .A2(_233_),
    .Z(_383_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _810_ (.I(_383_),
    .Z(_384_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _811_ (.A1(net13),
    .A2(_384_),
    .ZN(_385_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _812_ (.A1(\SPB[1] ),
    .A2(_381_),
    .ZN(_386_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _813_ (.A1(_385_),
    .A2(_386_),
    .B(_376_),
    .ZN(_061_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _814_ (.A1(_242_),
    .A2(_384_),
    .ZN(_387_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _815_ (.A1(_085_),
    .A2(_381_),
    .ZN(_388_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _816_ (.A1(_387_),
    .A2(_388_),
    .B(_376_),
    .ZN(_062_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _817_ (.A1(net15),
    .A2(_380_),
    .ZN(_389_));
 gf180mcu_fd_sc_mcu7t5v0__aoi211_1 _818_ (.A1(_087_),
    .A2(_381_),
    .B(_389_),
    .C(_147_),
    .ZN(_063_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _819_ (.A1(net16),
    .A2(_384_),
    .ZN(_390_));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 _820_ (.I(_380_),
    .Z(_391_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _821_ (.A1(\SPB[4] ),
    .A2(_391_),
    .ZN(_392_));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 _822_ (.I(_253_),
    .Z(_393_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _823_ (.A1(_390_),
    .A2(_392_),
    .B(_393_),
    .ZN(_064_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _824_ (.A1(net17),
    .A2(_384_),
    .ZN(_394_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _825_ (.A1(\SPB[5] ),
    .A2(_391_),
    .ZN(_395_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _826_ (.A1(_394_),
    .A2(_395_),
    .B(_393_),
    .ZN(_065_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _827_ (.A1(_218_),
    .A2(_383_),
    .ZN(_396_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _828_ (.A1(\SPB[6] ),
    .A2(_391_),
    .ZN(_397_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _829_ (.A1(_396_),
    .A2(_397_),
    .B(_393_),
    .ZN(_066_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _830_ (.A1(_223_),
    .A2(_383_),
    .ZN(_398_));
 gf180mcu_fd_sc_mcu7t5v0__nand2_1 _831_ (.A1(\SPB[7] ),
    .A2(_391_),
    .ZN(_399_));
 gf180mcu_fd_sc_mcu7t5v0__aoi21_1 _832_ (.A1(_398_),
    .A2(_399_),
    .B(_393_),
    .ZN(_067_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _833_ (.A1(_241_),
    .A2(_215_),
    .ZN(_068_));
 gf180mcu_fd_sc_mcu7t5v0__nor2_1 _834_ (.A1(_241_),
    .A2(_220_),
    .ZN(_069_));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _835_ (.D(_000_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(last_irq7_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _836_ (.D(_001_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net43));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _837_ (.D(_002_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net44));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _838_ (.D(_003_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(net45));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _839_ (.D(_004_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net46));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _840_ (.D(_005_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net47));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _841_ (.D(_006_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net48));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _842_ (.D(_007_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net49));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _843_ (.D(_008_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net50));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _844_ (.D(_009_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net83));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _845_ (.D(_010_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(net84));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _846_ (.D(_011_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(net85));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _847_ (.D(_012_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net86));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _848_ (.D(_013_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net87));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _849_ (.D(_014_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net88));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _850_ (.D(_015_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net89));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _851_ (.D(_016_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net90));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _852_ (.D(_017_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net91));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _853_ (.D(_018_),
    .CLK(clknet_3_4__leaf_wb_clk_i),
    .Q(net92));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _854_ (.D(_019_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(net93));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _855_ (.D(_020_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _856_ (.D(_021_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _857_ (.D(_022_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _858_ (.D(_023_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _859_ (.D(_024_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _860_ (.D(_025_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _861_ (.D(_026_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _862_ (.D(_027_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _863_ (.D(_028_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _864_ (.D(_029_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _865_ (.D(_030_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _866_ (.D(_031_),
    .CLK(clknet_3_0__leaf_wb_clk_i),
    .Q(\DDRB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _867_ (.D(_032_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _868_ (.D(_033_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _869_ (.D(_034_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\DDRB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _870_ (.D(_035_),
    .CLK(clknet_3_1__leaf_wb_clk_i),
    .Q(\DDRB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _871_ (.D(_036_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _872_ (.D(_037_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _873_ (.D(_038_),
    .CLK(clknet_3_5__leaf_wb_clk_i),
    .Q(\PORTA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _874_ (.D(_039_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _875_ (.D(_040_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _876_ (.D(_041_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _877_ (.D(_042_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _878_ (.D(_043_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _879_ (.D(_044_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _880_ (.D(_045_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _881_ (.D(_046_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _882_ (.D(_047_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _883_ (.D(_048_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\PORTB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _884_ (.D(_049_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _885_ (.D(_050_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _886_ (.D(_051_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\PORTB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _887_ (.D(_052_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\SPA[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _888_ (.D(_053_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPA[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _889_ (.D(_054_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(\SPA[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _890_ (.D(_055_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _891_ (.D(_056_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _892_ (.D(_057_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _893_ (.D(_058_),
    .CLK(clknet_3_2__leaf_wb_clk_i),
    .Q(\SPA[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _894_ (.D(_059_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\SPA[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _895_ (.D(_060_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(\SPB[0] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _896_ (.D(_061_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[1] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _897_ (.D(_062_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[2] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _898_ (.D(_063_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[3] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _899_ (.D(_064_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[4] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _900_ (.D(_065_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[5] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _901_ (.D(_066_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[6] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_2 _902_ (.D(_067_),
    .CLK(clknet_3_3__leaf_wb_clk_i),
    .Q(\SPB[7] ));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _903_ (.D(_068_),
    .CLK(clknet_3_7__leaf_wb_clk_i),
    .Q(last_irq0_trigger));
 gf180mcu_fd_sc_mcu7t5v0__dffq_1 _904_ (.D(_069_),
    .CLK(clknet_3_6__leaf_wb_clk_i),
    .Q(last_irg6_trigger));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_0_wb_clk_i (.I(wb_clk_i),
    .Z(clknet_0_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_0__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_0__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_1__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_1__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_2__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_2__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_3__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_3__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_4__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_4__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_5__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_5__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_6__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_6__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 clkbuf_3_7__f_wb_clk_i (.I(clknet_0_wb_clk_i),
    .Z(clknet_3_7__leaf_wb_clk_i));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold1 (.I(net92),
    .Z(net96));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold2 (.I(net87),
    .Z(net97));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold3 (.I(net89),
    .Z(net98));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold4 (.I(net86),
    .Z(net99));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold5 (.I(net88),
    .Z(net100));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold6 (.I(net93),
    .Z(net101));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 hold7 (.I(net90),
    .Z(net102));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 hold8 (.I(net91),
    .Z(net103));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input1 (.I(DAC_clk),
    .Z(net1));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input10 (.I(bus_cyc),
    .Z(net10));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input11 (.I(bus_we),
    .Z(net11));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input12 (.I(data_in[0]),
    .Z(net12));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input13 (.I(data_in[1]),
    .Z(net13));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input14 (.I(data_in[2]),
    .Z(net14));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input15 (.I(data_in[3]),
    .Z(net15));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input16 (.I(data_in[4]),
    .Z(net16));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input17 (.I(data_in[5]),
    .Z(net17));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input18 (.I(data_in[6]),
    .Z(net18));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input19 (.I(data_in[7]),
    .Z(net19));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input2 (.I(DAC_d1),
    .Z(net2));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input20 (.I(io_in[0]),
    .Z(net20));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input21 (.I(io_in[10]),
    .Z(net21));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input22 (.I(io_in[11]),
    .Z(net22));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input23 (.I(io_in[12]),
    .Z(net23));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input24 (.I(io_in[13]),
    .Z(net24));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input25 (.I(io_in[14]),
    .Z(net25));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input26 (.I(io_in[15]),
    .Z(net26));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input27 (.I(io_in[1]),
    .Z(net27));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input28 (.I(io_in[2]),
    .Z(net28));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input29 (.I(io_in[3]),
    .Z(net29));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input3 (.I(DAC_d2),
    .Z(net3));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input30 (.I(io_in[4]),
    .Z(net30));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input31 (.I(io_in[5]),
    .Z(net31));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input32 (.I(io_in[6]),
    .Z(net32));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input33 (.I(io_in[7]),
    .Z(net33));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input34 (.I(io_in[8]),
    .Z(net34));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input35 (.I(io_in[9]),
    .Z(net35));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input36 (.I(pwm0),
    .Z(net36));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input37 (.I(pwm1),
    .Z(net37));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input38 (.I(pwm2),
    .Z(net38));
 gf180mcu_fd_sc_mcu7t5v0__buf_2 input39 (.I(rst),
    .Z(net39));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input4 (.I(DAC_le),
    .Z(net4));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input40 (.I(tmr0_o),
    .Z(net40));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input41 (.I(tmr1_o),
    .Z(net41));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 input5 (.I(TXD),
    .Z(net5));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input6 (.I(addr[0]),
    .Z(net6));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input7 (.I(addr[1]),
    .Z(net7));
 gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 input8 (.I(addr[2]),
    .Z(net8));
 gf180mcu_fd_sc_mcu7t5v0__buf_1 input9 (.I(addr[3]),
    .Z(net9));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output42 (.I(net42),
    .Z(RXD));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output43 (.I(net43),
    .Z(data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output44 (.I(net44),
    .Z(data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output45 (.I(net45),
    .Z(data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output46 (.I(net46),
    .Z(data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output47 (.I(net47),
    .Z(data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output48 (.I(net48),
    .Z(data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output49 (.I(net49),
    .Z(data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output50 (.I(net50),
    .Z(data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output51 (.I(net51),
    .Z(io_oeb[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output52 (.I(net52),
    .Z(io_oeb[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output53 (.I(net53),
    .Z(io_oeb[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output54 (.I(net54),
    .Z(io_oeb[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output55 (.I(net55),
    .Z(io_oeb[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output56 (.I(net56),
    .Z(io_oeb[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output57 (.I(net57),
    .Z(io_oeb[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output58 (.I(net58),
    .Z(io_oeb[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output59 (.I(net59),
    .Z(io_oeb[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output60 (.I(net60),
    .Z(io_oeb[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output61 (.I(net61),
    .Z(io_oeb[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output62 (.I(net62),
    .Z(io_oeb[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output63 (.I(net63),
    .Z(io_oeb[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output64 (.I(net64),
    .Z(io_oeb[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output65 (.I(net65),
    .Z(io_oeb[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output66 (.I(net66),
    .Z(io_oeb[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output67 (.I(net67),
    .Z(io_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output68 (.I(net68),
    .Z(io_out[10]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output69 (.I(net69),
    .Z(io_out[11]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output70 (.I(net70),
    .Z(io_out[12]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output71 (.I(net71),
    .Z(io_out[13]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output72 (.I(net72),
    .Z(io_out[14]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output73 (.I(net73),
    .Z(io_out[15]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output74 (.I(net74),
    .Z(io_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output75 (.I(net75),
    .Z(io_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output76 (.I(net76),
    .Z(io_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output77 (.I(net77),
    .Z(io_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output78 (.I(net78),
    .Z(io_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output79 (.I(net79),
    .Z(io_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output80 (.I(net80),
    .Z(io_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output81 (.I(net81),
    .Z(io_out[8]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output82 (.I(net82),
    .Z(io_out[9]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output83 (.I(net83),
    .Z(irq0));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output84 (.I(net84),
    .Z(irq6));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output85 (.I(net85),
    .Z(irq7));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output86 (.I(net99),
    .Z(la_data_out[0]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output87 (.I(net97),
    .Z(la_data_out[1]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output88 (.I(net100),
    .Z(la_data_out[2]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output89 (.I(net98),
    .Z(la_data_out[3]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output90 (.I(net102),
    .Z(la_data_out[4]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output91 (.I(net103),
    .Z(la_data_out[5]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output92 (.I(net96),
    .Z(la_data_out[6]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output93 (.I(net101),
    .Z(la_data_out[7]));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output94 (.I(net94),
    .Z(tmr0_clk));
 gf180mcu_fd_sc_mcu7t5v0__buf_8 output95 (.I(net95),
    .Z(tmr1_clk));
endmodule

