magic
tech gf180mcuD
magscale 1 5
timestamp 1700750569
<< obsm1 >>
rect 672 1538 109312 73457
<< metal2 >>
rect 3472 74600 3528 75000
rect 5488 74600 5544 75000
rect 7504 74600 7560 75000
rect 9520 74600 9576 75000
rect 11536 74600 11592 75000
rect 13552 74600 13608 75000
rect 15568 74600 15624 75000
rect 17584 74600 17640 75000
rect 19600 74600 19656 75000
rect 21616 74600 21672 75000
rect 23632 74600 23688 75000
rect 25648 74600 25704 75000
rect 27664 74600 27720 75000
rect 29680 74600 29736 75000
rect 31696 74600 31752 75000
rect 33712 74600 33768 75000
rect 35728 74600 35784 75000
rect 37744 74600 37800 75000
rect 39760 74600 39816 75000
rect 41776 74600 41832 75000
rect 43792 74600 43848 75000
rect 45808 74600 45864 75000
rect 47824 74600 47880 75000
rect 49840 74600 49896 75000
rect 51856 74600 51912 75000
rect 53872 74600 53928 75000
rect 55888 74600 55944 75000
rect 57904 74600 57960 75000
rect 59920 74600 59976 75000
rect 61936 74600 61992 75000
rect 63952 74600 64008 75000
rect 65968 74600 66024 75000
rect 67984 74600 68040 75000
rect 70000 74600 70056 75000
rect 72016 74600 72072 75000
rect 74032 74600 74088 75000
rect 76048 74600 76104 75000
rect 78064 74600 78120 75000
rect 80080 74600 80136 75000
rect 82096 74600 82152 75000
rect 84112 74600 84168 75000
rect 86128 74600 86184 75000
rect 88144 74600 88200 75000
rect 90160 74600 90216 75000
rect 92176 74600 92232 75000
rect 94192 74600 94248 75000
rect 96208 74600 96264 75000
rect 98224 74600 98280 75000
rect 100240 74600 100296 75000
rect 102256 74600 102312 75000
rect 104272 74600 104328 75000
rect 106288 74600 106344 75000
rect 2464 0 2520 400
rect 3360 0 3416 400
rect 4256 0 4312 400
rect 5152 0 5208 400
rect 6048 0 6104 400
rect 6944 0 7000 400
rect 7840 0 7896 400
rect 8736 0 8792 400
rect 9632 0 9688 400
rect 10528 0 10584 400
rect 11424 0 11480 400
rect 12320 0 12376 400
rect 13216 0 13272 400
rect 14112 0 14168 400
rect 15008 0 15064 400
rect 15904 0 15960 400
rect 16800 0 16856 400
rect 17696 0 17752 400
rect 18592 0 18648 400
rect 19488 0 19544 400
rect 20384 0 20440 400
rect 21280 0 21336 400
rect 22176 0 22232 400
rect 23072 0 23128 400
rect 23968 0 24024 400
rect 24864 0 24920 400
rect 25760 0 25816 400
rect 26656 0 26712 400
rect 27552 0 27608 400
rect 28448 0 28504 400
rect 29344 0 29400 400
rect 30240 0 30296 400
rect 31136 0 31192 400
rect 32032 0 32088 400
rect 32928 0 32984 400
rect 33824 0 33880 400
rect 34720 0 34776 400
rect 35616 0 35672 400
rect 36512 0 36568 400
rect 37408 0 37464 400
rect 38304 0 38360 400
rect 39200 0 39256 400
rect 40096 0 40152 400
rect 40992 0 41048 400
rect 41888 0 41944 400
rect 42784 0 42840 400
rect 43680 0 43736 400
rect 44576 0 44632 400
rect 45472 0 45528 400
rect 46368 0 46424 400
rect 47264 0 47320 400
rect 48160 0 48216 400
rect 49056 0 49112 400
rect 49952 0 50008 400
rect 50848 0 50904 400
rect 51744 0 51800 400
rect 52640 0 52696 400
rect 53536 0 53592 400
rect 54432 0 54488 400
rect 55328 0 55384 400
rect 56224 0 56280 400
rect 57120 0 57176 400
rect 58016 0 58072 400
rect 58912 0 58968 400
rect 59808 0 59864 400
rect 60704 0 60760 400
rect 61600 0 61656 400
rect 62496 0 62552 400
rect 63392 0 63448 400
rect 64288 0 64344 400
rect 65184 0 65240 400
rect 66080 0 66136 400
rect 66976 0 67032 400
rect 67872 0 67928 400
rect 68768 0 68824 400
rect 69664 0 69720 400
rect 70560 0 70616 400
rect 71456 0 71512 400
rect 72352 0 72408 400
rect 73248 0 73304 400
rect 74144 0 74200 400
rect 75040 0 75096 400
rect 75936 0 75992 400
rect 76832 0 76888 400
rect 77728 0 77784 400
rect 78624 0 78680 400
rect 79520 0 79576 400
rect 80416 0 80472 400
rect 81312 0 81368 400
rect 82208 0 82264 400
rect 83104 0 83160 400
rect 84000 0 84056 400
rect 84896 0 84952 400
rect 85792 0 85848 400
rect 86688 0 86744 400
rect 87584 0 87640 400
rect 88480 0 88536 400
rect 89376 0 89432 400
rect 90272 0 90328 400
rect 91168 0 91224 400
rect 92064 0 92120 400
rect 92960 0 93016 400
rect 93856 0 93912 400
rect 94752 0 94808 400
rect 95648 0 95704 400
rect 96544 0 96600 400
rect 97440 0 97496 400
rect 98336 0 98392 400
rect 99232 0 99288 400
rect 100128 0 100184 400
rect 101024 0 101080 400
rect 101920 0 101976 400
rect 102816 0 102872 400
rect 103712 0 103768 400
rect 104608 0 104664 400
rect 105504 0 105560 400
rect 106400 0 106456 400
rect 107296 0 107352 400
<< obsm2 >>
rect 686 74570 3442 74600
rect 3558 74570 5458 74600
rect 5574 74570 7474 74600
rect 7590 74570 9490 74600
rect 9606 74570 11506 74600
rect 11622 74570 13522 74600
rect 13638 74570 15538 74600
rect 15654 74570 17554 74600
rect 17670 74570 19570 74600
rect 19686 74570 21586 74600
rect 21702 74570 23602 74600
rect 23718 74570 25618 74600
rect 25734 74570 27634 74600
rect 27750 74570 29650 74600
rect 29766 74570 31666 74600
rect 31782 74570 33682 74600
rect 33798 74570 35698 74600
rect 35814 74570 37714 74600
rect 37830 74570 39730 74600
rect 39846 74570 41746 74600
rect 41862 74570 43762 74600
rect 43878 74570 45778 74600
rect 45894 74570 47794 74600
rect 47910 74570 49810 74600
rect 49926 74570 51826 74600
rect 51942 74570 53842 74600
rect 53958 74570 55858 74600
rect 55974 74570 57874 74600
rect 57990 74570 59890 74600
rect 60006 74570 61906 74600
rect 62022 74570 63922 74600
rect 64038 74570 65938 74600
rect 66054 74570 67954 74600
rect 68070 74570 69970 74600
rect 70086 74570 71986 74600
rect 72102 74570 74002 74600
rect 74118 74570 76018 74600
rect 76134 74570 78034 74600
rect 78150 74570 80050 74600
rect 80166 74570 82066 74600
rect 82182 74570 84082 74600
rect 84198 74570 86098 74600
rect 86214 74570 88114 74600
rect 88230 74570 90130 74600
rect 90246 74570 92146 74600
rect 92262 74570 94162 74600
rect 94278 74570 96178 74600
rect 96294 74570 98194 74600
rect 98310 74570 100210 74600
rect 100326 74570 102226 74600
rect 102342 74570 104242 74600
rect 104358 74570 106258 74600
rect 106374 74570 109186 74600
rect 686 430 109186 74570
rect 686 350 2434 430
rect 2550 350 3330 430
rect 3446 350 4226 430
rect 4342 350 5122 430
rect 5238 350 6018 430
rect 6134 350 6914 430
rect 7030 350 7810 430
rect 7926 350 8706 430
rect 8822 350 9602 430
rect 9718 350 10498 430
rect 10614 350 11394 430
rect 11510 350 12290 430
rect 12406 350 13186 430
rect 13302 350 14082 430
rect 14198 350 14978 430
rect 15094 350 15874 430
rect 15990 350 16770 430
rect 16886 350 17666 430
rect 17782 350 18562 430
rect 18678 350 19458 430
rect 19574 350 20354 430
rect 20470 350 21250 430
rect 21366 350 22146 430
rect 22262 350 23042 430
rect 23158 350 23938 430
rect 24054 350 24834 430
rect 24950 350 25730 430
rect 25846 350 26626 430
rect 26742 350 27522 430
rect 27638 350 28418 430
rect 28534 350 29314 430
rect 29430 350 30210 430
rect 30326 350 31106 430
rect 31222 350 32002 430
rect 32118 350 32898 430
rect 33014 350 33794 430
rect 33910 350 34690 430
rect 34806 350 35586 430
rect 35702 350 36482 430
rect 36598 350 37378 430
rect 37494 350 38274 430
rect 38390 350 39170 430
rect 39286 350 40066 430
rect 40182 350 40962 430
rect 41078 350 41858 430
rect 41974 350 42754 430
rect 42870 350 43650 430
rect 43766 350 44546 430
rect 44662 350 45442 430
rect 45558 350 46338 430
rect 46454 350 47234 430
rect 47350 350 48130 430
rect 48246 350 49026 430
rect 49142 350 49922 430
rect 50038 350 50818 430
rect 50934 350 51714 430
rect 51830 350 52610 430
rect 52726 350 53506 430
rect 53622 350 54402 430
rect 54518 350 55298 430
rect 55414 350 56194 430
rect 56310 350 57090 430
rect 57206 350 57986 430
rect 58102 350 58882 430
rect 58998 350 59778 430
rect 59894 350 60674 430
rect 60790 350 61570 430
rect 61686 350 62466 430
rect 62582 350 63362 430
rect 63478 350 64258 430
rect 64374 350 65154 430
rect 65270 350 66050 430
rect 66166 350 66946 430
rect 67062 350 67842 430
rect 67958 350 68738 430
rect 68854 350 69634 430
rect 69750 350 70530 430
rect 70646 350 71426 430
rect 71542 350 72322 430
rect 72438 350 73218 430
rect 73334 350 74114 430
rect 74230 350 75010 430
rect 75126 350 75906 430
rect 76022 350 76802 430
rect 76918 350 77698 430
rect 77814 350 78594 430
rect 78710 350 79490 430
rect 79606 350 80386 430
rect 80502 350 81282 430
rect 81398 350 82178 430
rect 82294 350 83074 430
rect 83190 350 83970 430
rect 84086 350 84866 430
rect 84982 350 85762 430
rect 85878 350 86658 430
rect 86774 350 87554 430
rect 87670 350 88450 430
rect 88566 350 89346 430
rect 89462 350 90242 430
rect 90358 350 91138 430
rect 91254 350 92034 430
rect 92150 350 92930 430
rect 93046 350 93826 430
rect 93942 350 94722 430
rect 94838 350 95618 430
rect 95734 350 96514 430
rect 96630 350 97410 430
rect 97526 350 98306 430
rect 98422 350 99202 430
rect 99318 350 100098 430
rect 100214 350 100994 430
rect 101110 350 101890 430
rect 102006 350 102786 430
rect 102902 350 103682 430
rect 103798 350 104578 430
rect 104694 350 105474 430
rect 105590 350 106370 430
rect 106486 350 107266 430
rect 107382 350 109186 430
<< metal3 >>
rect 109600 72016 110000 72072
rect 109600 71344 110000 71400
rect 109600 70672 110000 70728
rect 0 70336 400 70392
rect 109600 70000 110000 70056
rect 0 69664 400 69720
rect 109600 69328 110000 69384
rect 0 68992 400 69048
rect 109600 68656 110000 68712
rect 0 68320 400 68376
rect 109600 67984 110000 68040
rect 0 67648 400 67704
rect 109600 67312 110000 67368
rect 0 66976 400 67032
rect 109600 66640 110000 66696
rect 0 66304 400 66360
rect 109600 65968 110000 66024
rect 0 65632 400 65688
rect 109600 65296 110000 65352
rect 0 64960 400 65016
rect 109600 64624 110000 64680
rect 0 64288 400 64344
rect 109600 63952 110000 64008
rect 0 63616 400 63672
rect 109600 63280 110000 63336
rect 0 62944 400 63000
rect 109600 62608 110000 62664
rect 0 62272 400 62328
rect 109600 61936 110000 61992
rect 0 61600 400 61656
rect 109600 61264 110000 61320
rect 0 60928 400 60984
rect 109600 60592 110000 60648
rect 0 60256 400 60312
rect 109600 59920 110000 59976
rect 0 59584 400 59640
rect 109600 59248 110000 59304
rect 0 58912 400 58968
rect 109600 58576 110000 58632
rect 0 58240 400 58296
rect 109600 57904 110000 57960
rect 0 57568 400 57624
rect 109600 57232 110000 57288
rect 0 56896 400 56952
rect 109600 56560 110000 56616
rect 0 56224 400 56280
rect 109600 55888 110000 55944
rect 0 55552 400 55608
rect 109600 55216 110000 55272
rect 0 54880 400 54936
rect 109600 54544 110000 54600
rect 0 54208 400 54264
rect 109600 53872 110000 53928
rect 0 53536 400 53592
rect 109600 53200 110000 53256
rect 0 52864 400 52920
rect 109600 52528 110000 52584
rect 0 52192 400 52248
rect 109600 51856 110000 51912
rect 0 51520 400 51576
rect 109600 51184 110000 51240
rect 0 50848 400 50904
rect 109600 50512 110000 50568
rect 0 50176 400 50232
rect 109600 49840 110000 49896
rect 0 49504 400 49560
rect 109600 49168 110000 49224
rect 0 48832 400 48888
rect 109600 48496 110000 48552
rect 0 48160 400 48216
rect 109600 47824 110000 47880
rect 0 47488 400 47544
rect 109600 47152 110000 47208
rect 0 46816 400 46872
rect 109600 46480 110000 46536
rect 0 46144 400 46200
rect 109600 45808 110000 45864
rect 0 45472 400 45528
rect 109600 45136 110000 45192
rect 0 44800 400 44856
rect 109600 44464 110000 44520
rect 0 44128 400 44184
rect 109600 43792 110000 43848
rect 0 43456 400 43512
rect 109600 43120 110000 43176
rect 0 42784 400 42840
rect 109600 42448 110000 42504
rect 0 42112 400 42168
rect 109600 41776 110000 41832
rect 0 41440 400 41496
rect 109600 41104 110000 41160
rect 0 40768 400 40824
rect 109600 40432 110000 40488
rect 0 40096 400 40152
rect 109600 39760 110000 39816
rect 0 39424 400 39480
rect 109600 39088 110000 39144
rect 0 38752 400 38808
rect 109600 38416 110000 38472
rect 0 38080 400 38136
rect 109600 37744 110000 37800
rect 0 37408 400 37464
rect 109600 37072 110000 37128
rect 0 36736 400 36792
rect 109600 36400 110000 36456
rect 0 36064 400 36120
rect 109600 35728 110000 35784
rect 0 35392 400 35448
rect 109600 35056 110000 35112
rect 0 34720 400 34776
rect 109600 34384 110000 34440
rect 0 34048 400 34104
rect 109600 33712 110000 33768
rect 0 33376 400 33432
rect 109600 33040 110000 33096
rect 0 32704 400 32760
rect 109600 32368 110000 32424
rect 0 32032 400 32088
rect 109600 31696 110000 31752
rect 0 31360 400 31416
rect 109600 31024 110000 31080
rect 0 30688 400 30744
rect 109600 30352 110000 30408
rect 0 30016 400 30072
rect 109600 29680 110000 29736
rect 0 29344 400 29400
rect 109600 29008 110000 29064
rect 0 28672 400 28728
rect 109600 28336 110000 28392
rect 0 28000 400 28056
rect 109600 27664 110000 27720
rect 0 27328 400 27384
rect 109600 26992 110000 27048
rect 0 26656 400 26712
rect 109600 26320 110000 26376
rect 0 25984 400 26040
rect 109600 25648 110000 25704
rect 0 25312 400 25368
rect 109600 24976 110000 25032
rect 0 24640 400 24696
rect 109600 24304 110000 24360
rect 0 23968 400 24024
rect 109600 23632 110000 23688
rect 0 23296 400 23352
rect 109600 22960 110000 23016
rect 0 22624 400 22680
rect 109600 22288 110000 22344
rect 0 21952 400 22008
rect 109600 21616 110000 21672
rect 0 21280 400 21336
rect 109600 20944 110000 21000
rect 0 20608 400 20664
rect 109600 20272 110000 20328
rect 0 19936 400 19992
rect 109600 19600 110000 19656
rect 0 19264 400 19320
rect 109600 18928 110000 18984
rect 0 18592 400 18648
rect 109600 18256 110000 18312
rect 0 17920 400 17976
rect 109600 17584 110000 17640
rect 0 17248 400 17304
rect 109600 16912 110000 16968
rect 0 16576 400 16632
rect 109600 16240 110000 16296
rect 0 15904 400 15960
rect 109600 15568 110000 15624
rect 0 15232 400 15288
rect 109600 14896 110000 14952
rect 0 14560 400 14616
rect 109600 14224 110000 14280
rect 0 13888 400 13944
rect 109600 13552 110000 13608
rect 0 13216 400 13272
rect 109600 12880 110000 12936
rect 0 12544 400 12600
rect 109600 12208 110000 12264
rect 0 11872 400 11928
rect 109600 11536 110000 11592
rect 0 11200 400 11256
rect 109600 10864 110000 10920
rect 0 10528 400 10584
rect 109600 10192 110000 10248
rect 0 9856 400 9912
rect 109600 9520 110000 9576
rect 0 9184 400 9240
rect 109600 8848 110000 8904
rect 0 8512 400 8568
rect 109600 8176 110000 8232
rect 0 7840 400 7896
rect 109600 7504 110000 7560
rect 0 7168 400 7224
rect 109600 6832 110000 6888
rect 0 6496 400 6552
rect 109600 6160 110000 6216
rect 0 5824 400 5880
rect 109600 5488 110000 5544
rect 0 5152 400 5208
rect 109600 4816 110000 4872
rect 0 4480 400 4536
rect 109600 4144 110000 4200
rect 109600 3472 110000 3528
rect 109600 2800 110000 2856
<< obsm3 >>
rect 400 72102 109634 73318
rect 400 71986 109570 72102
rect 400 71430 109634 71986
rect 400 71314 109570 71430
rect 400 70758 109634 71314
rect 400 70642 109570 70758
rect 400 70422 109634 70642
rect 430 70306 109634 70422
rect 400 70086 109634 70306
rect 400 69970 109570 70086
rect 400 69750 109634 69970
rect 430 69634 109634 69750
rect 400 69414 109634 69634
rect 400 69298 109570 69414
rect 400 69078 109634 69298
rect 430 68962 109634 69078
rect 400 68742 109634 68962
rect 400 68626 109570 68742
rect 400 68406 109634 68626
rect 430 68290 109634 68406
rect 400 68070 109634 68290
rect 400 67954 109570 68070
rect 400 67734 109634 67954
rect 430 67618 109634 67734
rect 400 67398 109634 67618
rect 400 67282 109570 67398
rect 400 67062 109634 67282
rect 430 66946 109634 67062
rect 400 66726 109634 66946
rect 400 66610 109570 66726
rect 400 66390 109634 66610
rect 430 66274 109634 66390
rect 400 66054 109634 66274
rect 400 65938 109570 66054
rect 400 65718 109634 65938
rect 430 65602 109634 65718
rect 400 65382 109634 65602
rect 400 65266 109570 65382
rect 400 65046 109634 65266
rect 430 64930 109634 65046
rect 400 64710 109634 64930
rect 400 64594 109570 64710
rect 400 64374 109634 64594
rect 430 64258 109634 64374
rect 400 64038 109634 64258
rect 400 63922 109570 64038
rect 400 63702 109634 63922
rect 430 63586 109634 63702
rect 400 63366 109634 63586
rect 400 63250 109570 63366
rect 400 63030 109634 63250
rect 430 62914 109634 63030
rect 400 62694 109634 62914
rect 400 62578 109570 62694
rect 400 62358 109634 62578
rect 430 62242 109634 62358
rect 400 62022 109634 62242
rect 400 61906 109570 62022
rect 400 61686 109634 61906
rect 430 61570 109634 61686
rect 400 61350 109634 61570
rect 400 61234 109570 61350
rect 400 61014 109634 61234
rect 430 60898 109634 61014
rect 400 60678 109634 60898
rect 400 60562 109570 60678
rect 400 60342 109634 60562
rect 430 60226 109634 60342
rect 400 60006 109634 60226
rect 400 59890 109570 60006
rect 400 59670 109634 59890
rect 430 59554 109634 59670
rect 400 59334 109634 59554
rect 400 59218 109570 59334
rect 400 58998 109634 59218
rect 430 58882 109634 58998
rect 400 58662 109634 58882
rect 400 58546 109570 58662
rect 400 58326 109634 58546
rect 430 58210 109634 58326
rect 400 57990 109634 58210
rect 400 57874 109570 57990
rect 400 57654 109634 57874
rect 430 57538 109634 57654
rect 400 57318 109634 57538
rect 400 57202 109570 57318
rect 400 56982 109634 57202
rect 430 56866 109634 56982
rect 400 56646 109634 56866
rect 400 56530 109570 56646
rect 400 56310 109634 56530
rect 430 56194 109634 56310
rect 400 55974 109634 56194
rect 400 55858 109570 55974
rect 400 55638 109634 55858
rect 430 55522 109634 55638
rect 400 55302 109634 55522
rect 400 55186 109570 55302
rect 400 54966 109634 55186
rect 430 54850 109634 54966
rect 400 54630 109634 54850
rect 400 54514 109570 54630
rect 400 54294 109634 54514
rect 430 54178 109634 54294
rect 400 53958 109634 54178
rect 400 53842 109570 53958
rect 400 53622 109634 53842
rect 430 53506 109634 53622
rect 400 53286 109634 53506
rect 400 53170 109570 53286
rect 400 52950 109634 53170
rect 430 52834 109634 52950
rect 400 52614 109634 52834
rect 400 52498 109570 52614
rect 400 52278 109634 52498
rect 430 52162 109634 52278
rect 400 51942 109634 52162
rect 400 51826 109570 51942
rect 400 51606 109634 51826
rect 430 51490 109634 51606
rect 400 51270 109634 51490
rect 400 51154 109570 51270
rect 400 50934 109634 51154
rect 430 50818 109634 50934
rect 400 50598 109634 50818
rect 400 50482 109570 50598
rect 400 50262 109634 50482
rect 430 50146 109634 50262
rect 400 49926 109634 50146
rect 400 49810 109570 49926
rect 400 49590 109634 49810
rect 430 49474 109634 49590
rect 400 49254 109634 49474
rect 400 49138 109570 49254
rect 400 48918 109634 49138
rect 430 48802 109634 48918
rect 400 48582 109634 48802
rect 400 48466 109570 48582
rect 400 48246 109634 48466
rect 430 48130 109634 48246
rect 400 47910 109634 48130
rect 400 47794 109570 47910
rect 400 47574 109634 47794
rect 430 47458 109634 47574
rect 400 47238 109634 47458
rect 400 47122 109570 47238
rect 400 46902 109634 47122
rect 430 46786 109634 46902
rect 400 46566 109634 46786
rect 400 46450 109570 46566
rect 400 46230 109634 46450
rect 430 46114 109634 46230
rect 400 45894 109634 46114
rect 400 45778 109570 45894
rect 400 45558 109634 45778
rect 430 45442 109634 45558
rect 400 45222 109634 45442
rect 400 45106 109570 45222
rect 400 44886 109634 45106
rect 430 44770 109634 44886
rect 400 44550 109634 44770
rect 400 44434 109570 44550
rect 400 44214 109634 44434
rect 430 44098 109634 44214
rect 400 43878 109634 44098
rect 400 43762 109570 43878
rect 400 43542 109634 43762
rect 430 43426 109634 43542
rect 400 43206 109634 43426
rect 400 43090 109570 43206
rect 400 42870 109634 43090
rect 430 42754 109634 42870
rect 400 42534 109634 42754
rect 400 42418 109570 42534
rect 400 42198 109634 42418
rect 430 42082 109634 42198
rect 400 41862 109634 42082
rect 400 41746 109570 41862
rect 400 41526 109634 41746
rect 430 41410 109634 41526
rect 400 41190 109634 41410
rect 400 41074 109570 41190
rect 400 40854 109634 41074
rect 430 40738 109634 40854
rect 400 40518 109634 40738
rect 400 40402 109570 40518
rect 400 40182 109634 40402
rect 430 40066 109634 40182
rect 400 39846 109634 40066
rect 400 39730 109570 39846
rect 400 39510 109634 39730
rect 430 39394 109634 39510
rect 400 39174 109634 39394
rect 400 39058 109570 39174
rect 400 38838 109634 39058
rect 430 38722 109634 38838
rect 400 38502 109634 38722
rect 400 38386 109570 38502
rect 400 38166 109634 38386
rect 430 38050 109634 38166
rect 400 37830 109634 38050
rect 400 37714 109570 37830
rect 400 37494 109634 37714
rect 430 37378 109634 37494
rect 400 37158 109634 37378
rect 400 37042 109570 37158
rect 400 36822 109634 37042
rect 430 36706 109634 36822
rect 400 36486 109634 36706
rect 400 36370 109570 36486
rect 400 36150 109634 36370
rect 430 36034 109634 36150
rect 400 35814 109634 36034
rect 400 35698 109570 35814
rect 400 35478 109634 35698
rect 430 35362 109634 35478
rect 400 35142 109634 35362
rect 400 35026 109570 35142
rect 400 34806 109634 35026
rect 430 34690 109634 34806
rect 400 34470 109634 34690
rect 400 34354 109570 34470
rect 400 34134 109634 34354
rect 430 34018 109634 34134
rect 400 33798 109634 34018
rect 400 33682 109570 33798
rect 400 33462 109634 33682
rect 430 33346 109634 33462
rect 400 33126 109634 33346
rect 400 33010 109570 33126
rect 400 32790 109634 33010
rect 430 32674 109634 32790
rect 400 32454 109634 32674
rect 400 32338 109570 32454
rect 400 32118 109634 32338
rect 430 32002 109634 32118
rect 400 31782 109634 32002
rect 400 31666 109570 31782
rect 400 31446 109634 31666
rect 430 31330 109634 31446
rect 400 31110 109634 31330
rect 400 30994 109570 31110
rect 400 30774 109634 30994
rect 430 30658 109634 30774
rect 400 30438 109634 30658
rect 400 30322 109570 30438
rect 400 30102 109634 30322
rect 430 29986 109634 30102
rect 400 29766 109634 29986
rect 400 29650 109570 29766
rect 400 29430 109634 29650
rect 430 29314 109634 29430
rect 400 29094 109634 29314
rect 400 28978 109570 29094
rect 400 28758 109634 28978
rect 430 28642 109634 28758
rect 400 28422 109634 28642
rect 400 28306 109570 28422
rect 400 28086 109634 28306
rect 430 27970 109634 28086
rect 400 27750 109634 27970
rect 400 27634 109570 27750
rect 400 27414 109634 27634
rect 430 27298 109634 27414
rect 400 27078 109634 27298
rect 400 26962 109570 27078
rect 400 26742 109634 26962
rect 430 26626 109634 26742
rect 400 26406 109634 26626
rect 400 26290 109570 26406
rect 400 26070 109634 26290
rect 430 25954 109634 26070
rect 400 25734 109634 25954
rect 400 25618 109570 25734
rect 400 25398 109634 25618
rect 430 25282 109634 25398
rect 400 25062 109634 25282
rect 400 24946 109570 25062
rect 400 24726 109634 24946
rect 430 24610 109634 24726
rect 400 24390 109634 24610
rect 400 24274 109570 24390
rect 400 24054 109634 24274
rect 430 23938 109634 24054
rect 400 23718 109634 23938
rect 400 23602 109570 23718
rect 400 23382 109634 23602
rect 430 23266 109634 23382
rect 400 23046 109634 23266
rect 400 22930 109570 23046
rect 400 22710 109634 22930
rect 430 22594 109634 22710
rect 400 22374 109634 22594
rect 400 22258 109570 22374
rect 400 22038 109634 22258
rect 430 21922 109634 22038
rect 400 21702 109634 21922
rect 400 21586 109570 21702
rect 400 21366 109634 21586
rect 430 21250 109634 21366
rect 400 21030 109634 21250
rect 400 20914 109570 21030
rect 400 20694 109634 20914
rect 430 20578 109634 20694
rect 400 20358 109634 20578
rect 400 20242 109570 20358
rect 400 20022 109634 20242
rect 430 19906 109634 20022
rect 400 19686 109634 19906
rect 400 19570 109570 19686
rect 400 19350 109634 19570
rect 430 19234 109634 19350
rect 400 19014 109634 19234
rect 400 18898 109570 19014
rect 400 18678 109634 18898
rect 430 18562 109634 18678
rect 400 18342 109634 18562
rect 400 18226 109570 18342
rect 400 18006 109634 18226
rect 430 17890 109634 18006
rect 400 17670 109634 17890
rect 400 17554 109570 17670
rect 400 17334 109634 17554
rect 430 17218 109634 17334
rect 400 16998 109634 17218
rect 400 16882 109570 16998
rect 400 16662 109634 16882
rect 430 16546 109634 16662
rect 400 16326 109634 16546
rect 400 16210 109570 16326
rect 400 15990 109634 16210
rect 430 15874 109634 15990
rect 400 15654 109634 15874
rect 400 15538 109570 15654
rect 400 15318 109634 15538
rect 430 15202 109634 15318
rect 400 14982 109634 15202
rect 400 14866 109570 14982
rect 400 14646 109634 14866
rect 430 14530 109634 14646
rect 400 14310 109634 14530
rect 400 14194 109570 14310
rect 400 13974 109634 14194
rect 430 13858 109634 13974
rect 400 13638 109634 13858
rect 400 13522 109570 13638
rect 400 13302 109634 13522
rect 430 13186 109634 13302
rect 400 12966 109634 13186
rect 400 12850 109570 12966
rect 400 12630 109634 12850
rect 430 12514 109634 12630
rect 400 12294 109634 12514
rect 400 12178 109570 12294
rect 400 11958 109634 12178
rect 430 11842 109634 11958
rect 400 11622 109634 11842
rect 400 11506 109570 11622
rect 400 11286 109634 11506
rect 430 11170 109634 11286
rect 400 10950 109634 11170
rect 400 10834 109570 10950
rect 400 10614 109634 10834
rect 430 10498 109634 10614
rect 400 10278 109634 10498
rect 400 10162 109570 10278
rect 400 9942 109634 10162
rect 430 9826 109634 9942
rect 400 9606 109634 9826
rect 400 9490 109570 9606
rect 400 9270 109634 9490
rect 430 9154 109634 9270
rect 400 8934 109634 9154
rect 400 8818 109570 8934
rect 400 8598 109634 8818
rect 430 8482 109634 8598
rect 400 8262 109634 8482
rect 400 8146 109570 8262
rect 400 7926 109634 8146
rect 430 7810 109634 7926
rect 400 7590 109634 7810
rect 400 7474 109570 7590
rect 400 7254 109634 7474
rect 430 7138 109634 7254
rect 400 6918 109634 7138
rect 400 6802 109570 6918
rect 400 6582 109634 6802
rect 430 6466 109634 6582
rect 400 6246 109634 6466
rect 400 6130 109570 6246
rect 400 5910 109634 6130
rect 430 5794 109634 5910
rect 400 5574 109634 5794
rect 400 5458 109570 5574
rect 400 5238 109634 5458
rect 430 5122 109634 5238
rect 400 4902 109634 5122
rect 400 4786 109570 4902
rect 400 4566 109634 4786
rect 430 4450 109634 4566
rect 400 4230 109634 4450
rect 400 4114 109570 4230
rect 400 3558 109634 4114
rect 400 3442 109570 3558
rect 400 2886 109634 3442
rect 400 2770 109570 2886
rect 400 1358 109634 2770
<< metal4 >>
rect 2224 1538 2384 73334
rect 9904 1538 10064 73334
rect 17584 1538 17744 73334
rect 25264 1538 25424 73334
rect 32944 1538 33104 73334
rect 40624 1538 40784 73334
rect 48304 1538 48464 73334
rect 55984 1538 56144 73334
rect 63664 1538 63824 73334
rect 71344 1538 71504 73334
rect 79024 1538 79184 73334
rect 86704 1538 86864 73334
rect 94384 1538 94544 73334
rect 102064 1538 102224 73334
<< obsm4 >>
rect 1862 1745 2194 64055
rect 2414 1745 9874 64055
rect 10094 1745 17554 64055
rect 17774 1745 25234 64055
rect 25454 1745 32914 64055
rect 33134 1745 40594 64055
rect 40814 1745 48274 64055
rect 48494 1745 55954 64055
rect 56174 1745 63634 64055
rect 63854 1745 71314 64055
rect 71534 1745 78994 64055
rect 79214 1745 86674 64055
rect 86894 1745 94354 64055
rect 94574 1745 102034 64055
rect 102254 1745 108178 64055
<< labels >>
rlabel metal3 s 0 43456 400 43512 6 RAM_end_addr[0]
port 1 nsew signal output
rlabel metal3 s 0 50176 400 50232 6 RAM_end_addr[10]
port 2 nsew signal output
rlabel metal3 s 0 50848 400 50904 6 RAM_end_addr[11]
port 3 nsew signal output
rlabel metal3 s 0 51520 400 51576 6 RAM_end_addr[12]
port 4 nsew signal output
rlabel metal3 s 0 52192 400 52248 6 RAM_end_addr[13]
port 5 nsew signal output
rlabel metal3 s 0 52864 400 52920 6 RAM_end_addr[14]
port 6 nsew signal output
rlabel metal3 s 0 53536 400 53592 6 RAM_end_addr[15]
port 7 nsew signal output
rlabel metal3 s 0 44128 400 44184 6 RAM_end_addr[1]
port 8 nsew signal output
rlabel metal3 s 0 44800 400 44856 6 RAM_end_addr[2]
port 9 nsew signal output
rlabel metal3 s 0 45472 400 45528 6 RAM_end_addr[3]
port 10 nsew signal output
rlabel metal3 s 0 46144 400 46200 6 RAM_end_addr[4]
port 11 nsew signal output
rlabel metal3 s 0 46816 400 46872 6 RAM_end_addr[5]
port 12 nsew signal output
rlabel metal3 s 0 47488 400 47544 6 RAM_end_addr[6]
port 13 nsew signal output
rlabel metal3 s 0 48160 400 48216 6 RAM_end_addr[7]
port 14 nsew signal output
rlabel metal3 s 0 48832 400 48888 6 RAM_end_addr[8]
port 15 nsew signal output
rlabel metal3 s 0 49504 400 49560 6 RAM_end_addr[9]
port 16 nsew signal output
rlabel metal3 s 0 30016 400 30072 6 RAM_start_addr[0]
port 17 nsew signal output
rlabel metal3 s 0 36736 400 36792 6 RAM_start_addr[10]
port 18 nsew signal output
rlabel metal3 s 0 37408 400 37464 6 RAM_start_addr[11]
port 19 nsew signal output
rlabel metal3 s 0 38080 400 38136 6 RAM_start_addr[12]
port 20 nsew signal output
rlabel metal3 s 0 38752 400 38808 6 RAM_start_addr[13]
port 21 nsew signal output
rlabel metal3 s 0 39424 400 39480 6 RAM_start_addr[14]
port 22 nsew signal output
rlabel metal3 s 0 40096 400 40152 6 RAM_start_addr[15]
port 23 nsew signal output
rlabel metal3 s 0 30688 400 30744 6 RAM_start_addr[1]
port 24 nsew signal output
rlabel metal3 s 0 31360 400 31416 6 RAM_start_addr[2]
port 25 nsew signal output
rlabel metal3 s 0 32032 400 32088 6 RAM_start_addr[3]
port 26 nsew signal output
rlabel metal3 s 0 32704 400 32760 6 RAM_start_addr[4]
port 27 nsew signal output
rlabel metal3 s 0 33376 400 33432 6 RAM_start_addr[5]
port 28 nsew signal output
rlabel metal3 s 0 34048 400 34104 6 RAM_start_addr[6]
port 29 nsew signal output
rlabel metal3 s 0 34720 400 34776 6 RAM_start_addr[7]
port 30 nsew signal output
rlabel metal3 s 0 35392 400 35448 6 RAM_start_addr[8]
port 31 nsew signal output
rlabel metal3 s 0 36064 400 36120 6 RAM_start_addr[9]
port 32 nsew signal output
rlabel metal2 s 102256 74600 102312 75000 6 WEb_raw
port 33 nsew signal output
rlabel metal3 s 0 42784 400 42840 6 boot_rom_en
port 34 nsew signal output
rlabel metal2 s 74032 74600 74088 75000 6 bus_addr[0]
port 35 nsew signal output
rlabel metal2 s 76048 74600 76104 75000 6 bus_addr[1]
port 36 nsew signal output
rlabel metal2 s 78064 74600 78120 75000 6 bus_addr[2]
port 37 nsew signal output
rlabel metal2 s 80080 74600 80136 75000 6 bus_addr[3]
port 38 nsew signal output
rlabel metal2 s 82096 74600 82152 75000 6 bus_addr[4]
port 39 nsew signal output
rlabel metal2 s 84112 74600 84168 75000 6 bus_addr[5]
port 40 nsew signal output
rlabel metal2 s 72016 74600 72072 75000 6 bus_cyc
port 41 nsew signal output
rlabel metal2 s 55888 74600 55944 75000 6 bus_data_out[0]
port 42 nsew signal output
rlabel metal2 s 57904 74600 57960 75000 6 bus_data_out[1]
port 43 nsew signal output
rlabel metal2 s 59920 74600 59976 75000 6 bus_data_out[2]
port 44 nsew signal output
rlabel metal2 s 61936 74600 61992 75000 6 bus_data_out[3]
port 45 nsew signal output
rlabel metal2 s 63952 74600 64008 75000 6 bus_data_out[4]
port 46 nsew signal output
rlabel metal2 s 65968 74600 66024 75000 6 bus_data_out[5]
port 47 nsew signal output
rlabel metal2 s 67984 74600 68040 75000 6 bus_data_out[6]
port 48 nsew signal output
rlabel metal2 s 70000 74600 70056 75000 6 bus_data_out[7]
port 49 nsew signal output
rlabel metal3 s 109600 43120 110000 43176 6 bus_in_gpios[0]
port 50 nsew signal input
rlabel metal3 s 109600 43792 110000 43848 6 bus_in_gpios[1]
port 51 nsew signal input
rlabel metal3 s 109600 44464 110000 44520 6 bus_in_gpios[2]
port 52 nsew signal input
rlabel metal3 s 109600 45136 110000 45192 6 bus_in_gpios[3]
port 53 nsew signal input
rlabel metal3 s 109600 45808 110000 45864 6 bus_in_gpios[4]
port 54 nsew signal input
rlabel metal3 s 109600 46480 110000 46536 6 bus_in_gpios[5]
port 55 nsew signal input
rlabel metal3 s 109600 47152 110000 47208 6 bus_in_gpios[6]
port 56 nsew signal input
rlabel metal3 s 109600 47824 110000 47880 6 bus_in_gpios[7]
port 57 nsew signal input
rlabel metal2 s 86128 74600 86184 75000 6 bus_in_serial_ports[0]
port 58 nsew signal input
rlabel metal2 s 88144 74600 88200 75000 6 bus_in_serial_ports[1]
port 59 nsew signal input
rlabel metal2 s 90160 74600 90216 75000 6 bus_in_serial_ports[2]
port 60 nsew signal input
rlabel metal2 s 92176 74600 92232 75000 6 bus_in_serial_ports[3]
port 61 nsew signal input
rlabel metal2 s 94192 74600 94248 75000 6 bus_in_serial_ports[4]
port 62 nsew signal input
rlabel metal2 s 96208 74600 96264 75000 6 bus_in_serial_ports[5]
port 63 nsew signal input
rlabel metal2 s 98224 74600 98280 75000 6 bus_in_serial_ports[6]
port 64 nsew signal input
rlabel metal2 s 100240 74600 100296 75000 6 bus_in_serial_ports[7]
port 65 nsew signal input
rlabel metal3 s 109600 56560 110000 56616 6 bus_in_sid[0]
port 66 nsew signal input
rlabel metal3 s 109600 57232 110000 57288 6 bus_in_sid[1]
port 67 nsew signal input
rlabel metal3 s 109600 57904 110000 57960 6 bus_in_sid[2]
port 68 nsew signal input
rlabel metal3 s 109600 58576 110000 58632 6 bus_in_sid[3]
port 69 nsew signal input
rlabel metal3 s 109600 59248 110000 59304 6 bus_in_sid[4]
port 70 nsew signal input
rlabel metal3 s 109600 59920 110000 59976 6 bus_in_sid[5]
port 71 nsew signal input
rlabel metal3 s 109600 60592 110000 60648 6 bus_in_sid[6]
port 72 nsew signal input
rlabel metal3 s 109600 61264 110000 61320 6 bus_in_sid[7]
port 73 nsew signal input
rlabel metal3 s 109600 50512 110000 50568 6 bus_in_timers[0]
port 74 nsew signal input
rlabel metal3 s 109600 51184 110000 51240 6 bus_in_timers[1]
port 75 nsew signal input
rlabel metal3 s 109600 51856 110000 51912 6 bus_in_timers[2]
port 76 nsew signal input
rlabel metal3 s 109600 52528 110000 52584 6 bus_in_timers[3]
port 77 nsew signal input
rlabel metal3 s 109600 53200 110000 53256 6 bus_in_timers[4]
port 78 nsew signal input
rlabel metal3 s 109600 53872 110000 53928 6 bus_in_timers[5]
port 79 nsew signal input
rlabel metal3 s 109600 54544 110000 54600 6 bus_in_timers[6]
port 80 nsew signal input
rlabel metal3 s 109600 55216 110000 55272 6 bus_in_timers[7]
port 81 nsew signal input
rlabel metal3 s 109600 42448 110000 42504 6 bus_we_gpios
port 82 nsew signal output
rlabel metal3 s 109600 49840 110000 49896 6 bus_we_serial_ports
port 83 nsew signal output
rlabel metal3 s 109600 55888 110000 55944 6 bus_we_sid
port 84 nsew signal output
rlabel metal3 s 109600 49168 110000 49224 6 bus_we_timers
port 85 nsew signal output
rlabel metal3 s 0 40768 400 40824 6 cs_port[0]
port 86 nsew signal output
rlabel metal3 s 0 41440 400 41496 6 cs_port[1]
port 87 nsew signal output
rlabel metal3 s 0 42112 400 42168 6 cs_port[2]
port 88 nsew signal output
rlabel metal2 s 3472 74600 3528 75000 6 io_in[0]
port 89 nsew signal input
rlabel metal2 s 23632 74600 23688 75000 6 io_in[10]
port 90 nsew signal input
rlabel metal2 s 25648 74600 25704 75000 6 io_in[11]
port 91 nsew signal input
rlabel metal2 s 27664 74600 27720 75000 6 io_in[12]
port 92 nsew signal input
rlabel metal2 s 29680 74600 29736 75000 6 io_in[13]
port 93 nsew signal input
rlabel metal2 s 31696 74600 31752 75000 6 io_in[14]
port 94 nsew signal input
rlabel metal2 s 33712 74600 33768 75000 6 io_in[15]
port 95 nsew signal input
rlabel metal2 s 35728 74600 35784 75000 6 io_in[16]
port 96 nsew signal input
rlabel metal2 s 37744 74600 37800 75000 6 io_in[17]
port 97 nsew signal input
rlabel metal2 s 39760 74600 39816 75000 6 io_in[18]
port 98 nsew signal input
rlabel metal2 s 5488 74600 5544 75000 6 io_in[1]
port 99 nsew signal input
rlabel metal2 s 7504 74600 7560 75000 6 io_in[2]
port 100 nsew signal input
rlabel metal2 s 9520 74600 9576 75000 6 io_in[3]
port 101 nsew signal input
rlabel metal2 s 11536 74600 11592 75000 6 io_in[4]
port 102 nsew signal input
rlabel metal2 s 13552 74600 13608 75000 6 io_in[5]
port 103 nsew signal input
rlabel metal2 s 15568 74600 15624 75000 6 io_in[6]
port 104 nsew signal input
rlabel metal2 s 17584 74600 17640 75000 6 io_in[7]
port 105 nsew signal input
rlabel metal2 s 19600 74600 19656 75000 6 io_in[8]
port 106 nsew signal input
rlabel metal2 s 21616 74600 21672 75000 6 io_in[9]
port 107 nsew signal input
rlabel metal3 s 0 17248 400 17304 6 io_oeb[0]
port 108 nsew signal output
rlabel metal3 s 0 23968 400 24024 6 io_oeb[10]
port 109 nsew signal output
rlabel metal3 s 0 24640 400 24696 6 io_oeb[11]
port 110 nsew signal output
rlabel metal3 s 0 25312 400 25368 6 io_oeb[12]
port 111 nsew signal output
rlabel metal3 s 0 25984 400 26040 6 io_oeb[13]
port 112 nsew signal output
rlabel metal3 s 0 26656 400 26712 6 io_oeb[14]
port 113 nsew signal output
rlabel metal3 s 0 27328 400 27384 6 io_oeb[15]
port 114 nsew signal output
rlabel metal3 s 0 28000 400 28056 6 io_oeb[16]
port 115 nsew signal output
rlabel metal3 s 0 28672 400 28728 6 io_oeb[17]
port 116 nsew signal output
rlabel metal3 s 0 29344 400 29400 6 io_oeb[18]
port 117 nsew signal output
rlabel metal3 s 0 17920 400 17976 6 io_oeb[1]
port 118 nsew signal output
rlabel metal3 s 0 18592 400 18648 6 io_oeb[2]
port 119 nsew signal output
rlabel metal3 s 0 19264 400 19320 6 io_oeb[3]
port 120 nsew signal output
rlabel metal3 s 0 19936 400 19992 6 io_oeb[4]
port 121 nsew signal output
rlabel metal3 s 0 20608 400 20664 6 io_oeb[5]
port 122 nsew signal output
rlabel metal3 s 0 21280 400 21336 6 io_oeb[6]
port 123 nsew signal output
rlabel metal3 s 0 21952 400 22008 6 io_oeb[7]
port 124 nsew signal output
rlabel metal3 s 0 22624 400 22680 6 io_oeb[8]
port 125 nsew signal output
rlabel metal3 s 0 23296 400 23352 6 io_oeb[9]
port 126 nsew signal output
rlabel metal3 s 0 4480 400 4536 6 io_out[0]
port 127 nsew signal output
rlabel metal3 s 0 11200 400 11256 6 io_out[10]
port 128 nsew signal output
rlabel metal3 s 0 11872 400 11928 6 io_out[11]
port 129 nsew signal output
rlabel metal3 s 0 12544 400 12600 6 io_out[12]
port 130 nsew signal output
rlabel metal3 s 0 13216 400 13272 6 io_out[13]
port 131 nsew signal output
rlabel metal3 s 0 13888 400 13944 6 io_out[14]
port 132 nsew signal output
rlabel metal3 s 0 14560 400 14616 6 io_out[15]
port 133 nsew signal output
rlabel metal3 s 0 15232 400 15288 6 io_out[16]
port 134 nsew signal output
rlabel metal3 s 0 15904 400 15960 6 io_out[17]
port 135 nsew signal output
rlabel metal3 s 0 16576 400 16632 6 io_out[18]
port 136 nsew signal output
rlabel metal3 s 0 5152 400 5208 6 io_out[1]
port 137 nsew signal output
rlabel metal3 s 0 5824 400 5880 6 io_out[2]
port 138 nsew signal output
rlabel metal3 s 0 6496 400 6552 6 io_out[3]
port 139 nsew signal output
rlabel metal3 s 0 7168 400 7224 6 io_out[4]
port 140 nsew signal output
rlabel metal3 s 0 7840 400 7896 6 io_out[5]
port 141 nsew signal output
rlabel metal3 s 0 8512 400 8568 6 io_out[6]
port 142 nsew signal output
rlabel metal3 s 0 9184 400 9240 6 io_out[7]
port 143 nsew signal output
rlabel metal3 s 0 9856 400 9912 6 io_out[8]
port 144 nsew signal output
rlabel metal3 s 0 10528 400 10584 6 io_out[9]
port 145 nsew signal output
rlabel metal3 s 109600 40432 110000 40488 6 irq[0]
port 146 nsew signal output
rlabel metal3 s 109600 41104 110000 41160 6 irq[1]
port 147 nsew signal output
rlabel metal3 s 109600 41776 110000 41832 6 irq[2]
port 148 nsew signal output
rlabel metal2 s 41776 74600 41832 75000 6 irqs[0]
port 149 nsew signal input
rlabel metal2 s 43792 74600 43848 75000 6 irqs[1]
port 150 nsew signal input
rlabel metal2 s 45808 74600 45864 75000 6 irqs[2]
port 151 nsew signal input
rlabel metal2 s 47824 74600 47880 75000 6 irqs[3]
port 152 nsew signal input
rlabel metal2 s 49840 74600 49896 75000 6 irqs[4]
port 153 nsew signal input
rlabel metal2 s 51856 74600 51912 75000 6 irqs[5]
port 154 nsew signal input
rlabel metal2 s 53872 74600 53928 75000 6 irqs[6]
port 155 nsew signal input
rlabel metal3 s 109600 2800 110000 2856 6 la_data_out[0]
port 156 nsew signal output
rlabel metal3 s 109600 9520 110000 9576 6 la_data_out[10]
port 157 nsew signal output
rlabel metal3 s 109600 10192 110000 10248 6 la_data_out[11]
port 158 nsew signal output
rlabel metal3 s 109600 10864 110000 10920 6 la_data_out[12]
port 159 nsew signal output
rlabel metal3 s 109600 11536 110000 11592 6 la_data_out[13]
port 160 nsew signal output
rlabel metal3 s 109600 12208 110000 12264 6 la_data_out[14]
port 161 nsew signal output
rlabel metal3 s 109600 12880 110000 12936 6 la_data_out[15]
port 162 nsew signal output
rlabel metal3 s 109600 13552 110000 13608 6 la_data_out[16]
port 163 nsew signal output
rlabel metal3 s 109600 14224 110000 14280 6 la_data_out[17]
port 164 nsew signal output
rlabel metal3 s 109600 14896 110000 14952 6 la_data_out[18]
port 165 nsew signal output
rlabel metal3 s 109600 15568 110000 15624 6 la_data_out[19]
port 166 nsew signal output
rlabel metal3 s 109600 3472 110000 3528 6 la_data_out[1]
port 167 nsew signal output
rlabel metal3 s 109600 16240 110000 16296 6 la_data_out[20]
port 168 nsew signal output
rlabel metal3 s 109600 16912 110000 16968 6 la_data_out[21]
port 169 nsew signal output
rlabel metal3 s 109600 17584 110000 17640 6 la_data_out[22]
port 170 nsew signal output
rlabel metal3 s 109600 18256 110000 18312 6 la_data_out[23]
port 171 nsew signal output
rlabel metal3 s 109600 18928 110000 18984 6 la_data_out[24]
port 172 nsew signal output
rlabel metal3 s 109600 19600 110000 19656 6 la_data_out[25]
port 173 nsew signal output
rlabel metal3 s 109600 20272 110000 20328 6 la_data_out[26]
port 174 nsew signal output
rlabel metal3 s 109600 20944 110000 21000 6 la_data_out[27]
port 175 nsew signal output
rlabel metal3 s 109600 21616 110000 21672 6 la_data_out[28]
port 176 nsew signal output
rlabel metal3 s 109600 22288 110000 22344 6 la_data_out[29]
port 177 nsew signal output
rlabel metal3 s 109600 4144 110000 4200 6 la_data_out[2]
port 178 nsew signal output
rlabel metal3 s 109600 22960 110000 23016 6 la_data_out[30]
port 179 nsew signal output
rlabel metal3 s 109600 23632 110000 23688 6 la_data_out[31]
port 180 nsew signal output
rlabel metal3 s 109600 24304 110000 24360 6 la_data_out[32]
port 181 nsew signal output
rlabel metal3 s 109600 24976 110000 25032 6 la_data_out[33]
port 182 nsew signal output
rlabel metal3 s 109600 25648 110000 25704 6 la_data_out[34]
port 183 nsew signal output
rlabel metal3 s 109600 26320 110000 26376 6 la_data_out[35]
port 184 nsew signal output
rlabel metal3 s 109600 26992 110000 27048 6 la_data_out[36]
port 185 nsew signal output
rlabel metal3 s 109600 27664 110000 27720 6 la_data_out[37]
port 186 nsew signal output
rlabel metal3 s 109600 28336 110000 28392 6 la_data_out[38]
port 187 nsew signal output
rlabel metal3 s 109600 29008 110000 29064 6 la_data_out[39]
port 188 nsew signal output
rlabel metal3 s 109600 4816 110000 4872 6 la_data_out[3]
port 189 nsew signal output
rlabel metal3 s 109600 29680 110000 29736 6 la_data_out[40]
port 190 nsew signal output
rlabel metal3 s 109600 30352 110000 30408 6 la_data_out[41]
port 191 nsew signal output
rlabel metal3 s 109600 31024 110000 31080 6 la_data_out[42]
port 192 nsew signal output
rlabel metal3 s 109600 31696 110000 31752 6 la_data_out[43]
port 193 nsew signal output
rlabel metal3 s 109600 32368 110000 32424 6 la_data_out[44]
port 194 nsew signal output
rlabel metal3 s 109600 33040 110000 33096 6 la_data_out[45]
port 195 nsew signal output
rlabel metal3 s 109600 33712 110000 33768 6 la_data_out[46]
port 196 nsew signal output
rlabel metal3 s 109600 34384 110000 34440 6 la_data_out[47]
port 197 nsew signal output
rlabel metal3 s 109600 35056 110000 35112 6 la_data_out[48]
port 198 nsew signal output
rlabel metal3 s 109600 35728 110000 35784 6 la_data_out[49]
port 199 nsew signal output
rlabel metal3 s 109600 5488 110000 5544 6 la_data_out[4]
port 200 nsew signal output
rlabel metal3 s 109600 36400 110000 36456 6 la_data_out[50]
port 201 nsew signal output
rlabel metal3 s 109600 37072 110000 37128 6 la_data_out[51]
port 202 nsew signal output
rlabel metal3 s 109600 37744 110000 37800 6 la_data_out[52]
port 203 nsew signal output
rlabel metal3 s 109600 38416 110000 38472 6 la_data_out[53]
port 204 nsew signal output
rlabel metal3 s 109600 39088 110000 39144 6 la_data_out[54]
port 205 nsew signal output
rlabel metal3 s 109600 39760 110000 39816 6 la_data_out[55]
port 206 nsew signal output
rlabel metal3 s 109600 6160 110000 6216 6 la_data_out[5]
port 207 nsew signal output
rlabel metal3 s 109600 6832 110000 6888 6 la_data_out[6]
port 208 nsew signal output
rlabel metal3 s 109600 7504 110000 7560 6 la_data_out[7]
port 209 nsew signal output
rlabel metal3 s 109600 8176 110000 8232 6 la_data_out[8]
port 210 nsew signal output
rlabel metal3 s 109600 8848 110000 8904 6 la_data_out[9]
port 211 nsew signal output
rlabel metal2 s 93856 0 93912 400 6 last_addr[0]
port 212 nsew signal output
rlabel metal2 s 102816 0 102872 400 6 last_addr[10]
port 213 nsew signal output
rlabel metal2 s 103712 0 103768 400 6 last_addr[11]
port 214 nsew signal output
rlabel metal2 s 104608 0 104664 400 6 last_addr[12]
port 215 nsew signal output
rlabel metal2 s 105504 0 105560 400 6 last_addr[13]
port 216 nsew signal output
rlabel metal2 s 106400 0 106456 400 6 last_addr[14]
port 217 nsew signal output
rlabel metal2 s 107296 0 107352 400 6 last_addr[15]
port 218 nsew signal output
rlabel metal2 s 94752 0 94808 400 6 last_addr[1]
port 219 nsew signal output
rlabel metal2 s 95648 0 95704 400 6 last_addr[2]
port 220 nsew signal output
rlabel metal2 s 96544 0 96600 400 6 last_addr[3]
port 221 nsew signal output
rlabel metal2 s 97440 0 97496 400 6 last_addr[4]
port 222 nsew signal output
rlabel metal2 s 98336 0 98392 400 6 last_addr[5]
port 223 nsew signal output
rlabel metal2 s 99232 0 99288 400 6 last_addr[6]
port 224 nsew signal output
rlabel metal2 s 100128 0 100184 400 6 last_addr[7]
port 225 nsew signal output
rlabel metal2 s 101024 0 101080 400 6 last_addr[8]
port 226 nsew signal output
rlabel metal2 s 101920 0 101976 400 6 last_addr[9]
port 227 nsew signal output
rlabel metal2 s 106288 74600 106344 75000 6 le_hi_act
port 228 nsew signal output
rlabel metal2 s 104272 74600 104328 75000 6 le_lo_act
port 229 nsew signal output
rlabel metal3 s 0 64960 400 65016 6 ram_bus_in[0]
port 230 nsew signal input
rlabel metal3 s 0 65632 400 65688 6 ram_bus_in[1]
port 231 nsew signal input
rlabel metal3 s 0 66304 400 66360 6 ram_bus_in[2]
port 232 nsew signal input
rlabel metal3 s 0 66976 400 67032 6 ram_bus_in[3]
port 233 nsew signal input
rlabel metal3 s 0 67648 400 67704 6 ram_bus_in[4]
port 234 nsew signal input
rlabel metal3 s 0 68320 400 68376 6 ram_bus_in[5]
port 235 nsew signal input
rlabel metal3 s 0 68992 400 69048 6 ram_bus_in[6]
port 236 nsew signal input
rlabel metal3 s 0 69664 400 69720 6 ram_bus_in[7]
port 237 nsew signal input
rlabel metal3 s 0 70336 400 70392 6 ram_enabled
port 238 nsew signal output
rlabel metal3 s 109600 61936 110000 61992 6 requested_addr[0]
port 239 nsew signal output
rlabel metal3 s 109600 68656 110000 68712 6 requested_addr[10]
port 240 nsew signal output
rlabel metal3 s 109600 69328 110000 69384 6 requested_addr[11]
port 241 nsew signal output
rlabel metal3 s 109600 70000 110000 70056 6 requested_addr[12]
port 242 nsew signal output
rlabel metal3 s 109600 70672 110000 70728 6 requested_addr[13]
port 243 nsew signal output
rlabel metal3 s 109600 71344 110000 71400 6 requested_addr[14]
port 244 nsew signal output
rlabel metal3 s 109600 72016 110000 72072 6 requested_addr[15]
port 245 nsew signal output
rlabel metal3 s 109600 62608 110000 62664 6 requested_addr[1]
port 246 nsew signal output
rlabel metal3 s 109600 63280 110000 63336 6 requested_addr[2]
port 247 nsew signal output
rlabel metal3 s 109600 63952 110000 64008 6 requested_addr[3]
port 248 nsew signal output
rlabel metal3 s 109600 64624 110000 64680 6 requested_addr[4]
port 249 nsew signal output
rlabel metal3 s 109600 65296 110000 65352 6 requested_addr[5]
port 250 nsew signal output
rlabel metal3 s 109600 65968 110000 66024 6 requested_addr[6]
port 251 nsew signal output
rlabel metal3 s 109600 66640 110000 66696 6 requested_addr[7]
port 252 nsew signal output
rlabel metal3 s 109600 67312 110000 67368 6 requested_addr[8]
port 253 nsew signal output
rlabel metal3 s 109600 67984 110000 68040 6 requested_addr[9]
port 254 nsew signal output
rlabel metal3 s 109600 48496 110000 48552 6 reset_out
port 255 nsew signal output
rlabel metal3 s 0 59584 400 59640 6 rom_bus_in[0]
port 256 nsew signal input
rlabel metal3 s 0 60256 400 60312 6 rom_bus_in[1]
port 257 nsew signal input
rlabel metal3 s 0 60928 400 60984 6 rom_bus_in[2]
port 258 nsew signal input
rlabel metal3 s 0 61600 400 61656 6 rom_bus_in[3]
port 259 nsew signal input
rlabel metal3 s 0 62272 400 62328 6 rom_bus_in[4]
port 260 nsew signal input
rlabel metal3 s 0 62944 400 63000 6 rom_bus_in[5]
port 261 nsew signal input
rlabel metal3 s 0 63616 400 63672 6 rom_bus_in[6]
port 262 nsew signal input
rlabel metal3 s 0 64288 400 64344 6 rom_bus_in[7]
port 263 nsew signal input
rlabel metal3 s 0 54208 400 54264 6 rom_bus_out[0]
port 264 nsew signal output
rlabel metal3 s 0 54880 400 54936 6 rom_bus_out[1]
port 265 nsew signal output
rlabel metal3 s 0 55552 400 55608 6 rom_bus_out[2]
port 266 nsew signal output
rlabel metal3 s 0 56224 400 56280 6 rom_bus_out[3]
port 267 nsew signal output
rlabel metal3 s 0 56896 400 56952 6 rom_bus_out[4]
port 268 nsew signal output
rlabel metal3 s 0 57568 400 57624 6 rom_bus_out[5]
port 269 nsew signal output
rlabel metal3 s 0 58240 400 58296 6 rom_bus_out[6]
port 270 nsew signal output
rlabel metal3 s 0 58912 400 58968 6 rom_bus_out[7]
port 271 nsew signal output
rlabel metal4 s 2224 1538 2384 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 32944 1538 33104 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 48304 1538 48464 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 63664 1538 63824 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 79024 1538 79184 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 94384 1538 94544 73334 6 vdd
port 272 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 25264 1538 25424 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 40624 1538 40784 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 55984 1538 56144 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 71344 1538 71504 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 86704 1538 86864 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal4 s 102064 1538 102224 73334 6 vss
port 273 nsew ground bidirectional
rlabel metal2 s 2464 0 2520 400 6 wb_clk_i
port 274 nsew signal input
rlabel metal2 s 3360 0 3416 400 6 wb_rst_i
port 275 nsew signal input
rlabel metal2 s 4256 0 4312 400 6 wbs_ack_o
port 276 nsew signal output
rlabel metal2 s 7840 0 7896 400 6 wbs_adr_i[0]
port 277 nsew signal input
rlabel metal2 s 34720 0 34776 400 6 wbs_adr_i[10]
port 278 nsew signal input
rlabel metal2 s 37408 0 37464 400 6 wbs_adr_i[11]
port 279 nsew signal input
rlabel metal2 s 40096 0 40152 400 6 wbs_adr_i[12]
port 280 nsew signal input
rlabel metal2 s 42784 0 42840 400 6 wbs_adr_i[13]
port 281 nsew signal input
rlabel metal2 s 45472 0 45528 400 6 wbs_adr_i[14]
port 282 nsew signal input
rlabel metal2 s 48160 0 48216 400 6 wbs_adr_i[15]
port 283 nsew signal input
rlabel metal2 s 50848 0 50904 400 6 wbs_adr_i[16]
port 284 nsew signal input
rlabel metal2 s 53536 0 53592 400 6 wbs_adr_i[17]
port 285 nsew signal input
rlabel metal2 s 56224 0 56280 400 6 wbs_adr_i[18]
port 286 nsew signal input
rlabel metal2 s 58912 0 58968 400 6 wbs_adr_i[19]
port 287 nsew signal input
rlabel metal2 s 10528 0 10584 400 6 wbs_adr_i[1]
port 288 nsew signal input
rlabel metal2 s 61600 0 61656 400 6 wbs_adr_i[20]
port 289 nsew signal input
rlabel metal2 s 64288 0 64344 400 6 wbs_adr_i[21]
port 290 nsew signal input
rlabel metal2 s 66976 0 67032 400 6 wbs_adr_i[22]
port 291 nsew signal input
rlabel metal2 s 69664 0 69720 400 6 wbs_adr_i[23]
port 292 nsew signal input
rlabel metal2 s 72352 0 72408 400 6 wbs_adr_i[24]
port 293 nsew signal input
rlabel metal2 s 75040 0 75096 400 6 wbs_adr_i[25]
port 294 nsew signal input
rlabel metal2 s 77728 0 77784 400 6 wbs_adr_i[26]
port 295 nsew signal input
rlabel metal2 s 80416 0 80472 400 6 wbs_adr_i[27]
port 296 nsew signal input
rlabel metal2 s 83104 0 83160 400 6 wbs_adr_i[28]
port 297 nsew signal input
rlabel metal2 s 85792 0 85848 400 6 wbs_adr_i[29]
port 298 nsew signal input
rlabel metal2 s 13216 0 13272 400 6 wbs_adr_i[2]
port 299 nsew signal input
rlabel metal2 s 88480 0 88536 400 6 wbs_adr_i[30]
port 300 nsew signal input
rlabel metal2 s 91168 0 91224 400 6 wbs_adr_i[31]
port 301 nsew signal input
rlabel metal2 s 15904 0 15960 400 6 wbs_adr_i[3]
port 302 nsew signal input
rlabel metal2 s 18592 0 18648 400 6 wbs_adr_i[4]
port 303 nsew signal input
rlabel metal2 s 21280 0 21336 400 6 wbs_adr_i[5]
port 304 nsew signal input
rlabel metal2 s 23968 0 24024 400 6 wbs_adr_i[6]
port 305 nsew signal input
rlabel metal2 s 26656 0 26712 400 6 wbs_adr_i[7]
port 306 nsew signal input
rlabel metal2 s 29344 0 29400 400 6 wbs_adr_i[8]
port 307 nsew signal input
rlabel metal2 s 32032 0 32088 400 6 wbs_adr_i[9]
port 308 nsew signal input
rlabel metal2 s 5152 0 5208 400 6 wbs_cyc_i
port 309 nsew signal input
rlabel metal2 s 8736 0 8792 400 6 wbs_dat_i[0]
port 310 nsew signal input
rlabel metal2 s 35616 0 35672 400 6 wbs_dat_i[10]
port 311 nsew signal input
rlabel metal2 s 38304 0 38360 400 6 wbs_dat_i[11]
port 312 nsew signal input
rlabel metal2 s 40992 0 41048 400 6 wbs_dat_i[12]
port 313 nsew signal input
rlabel metal2 s 43680 0 43736 400 6 wbs_dat_i[13]
port 314 nsew signal input
rlabel metal2 s 46368 0 46424 400 6 wbs_dat_i[14]
port 315 nsew signal input
rlabel metal2 s 49056 0 49112 400 6 wbs_dat_i[15]
port 316 nsew signal input
rlabel metal2 s 51744 0 51800 400 6 wbs_dat_i[16]
port 317 nsew signal input
rlabel metal2 s 54432 0 54488 400 6 wbs_dat_i[17]
port 318 nsew signal input
rlabel metal2 s 57120 0 57176 400 6 wbs_dat_i[18]
port 319 nsew signal input
rlabel metal2 s 59808 0 59864 400 6 wbs_dat_i[19]
port 320 nsew signal input
rlabel metal2 s 11424 0 11480 400 6 wbs_dat_i[1]
port 321 nsew signal input
rlabel metal2 s 62496 0 62552 400 6 wbs_dat_i[20]
port 322 nsew signal input
rlabel metal2 s 65184 0 65240 400 6 wbs_dat_i[21]
port 323 nsew signal input
rlabel metal2 s 67872 0 67928 400 6 wbs_dat_i[22]
port 324 nsew signal input
rlabel metal2 s 70560 0 70616 400 6 wbs_dat_i[23]
port 325 nsew signal input
rlabel metal2 s 73248 0 73304 400 6 wbs_dat_i[24]
port 326 nsew signal input
rlabel metal2 s 75936 0 75992 400 6 wbs_dat_i[25]
port 327 nsew signal input
rlabel metal2 s 78624 0 78680 400 6 wbs_dat_i[26]
port 328 nsew signal input
rlabel metal2 s 81312 0 81368 400 6 wbs_dat_i[27]
port 329 nsew signal input
rlabel metal2 s 84000 0 84056 400 6 wbs_dat_i[28]
port 330 nsew signal input
rlabel metal2 s 86688 0 86744 400 6 wbs_dat_i[29]
port 331 nsew signal input
rlabel metal2 s 14112 0 14168 400 6 wbs_dat_i[2]
port 332 nsew signal input
rlabel metal2 s 89376 0 89432 400 6 wbs_dat_i[30]
port 333 nsew signal input
rlabel metal2 s 92064 0 92120 400 6 wbs_dat_i[31]
port 334 nsew signal input
rlabel metal2 s 16800 0 16856 400 6 wbs_dat_i[3]
port 335 nsew signal input
rlabel metal2 s 19488 0 19544 400 6 wbs_dat_i[4]
port 336 nsew signal input
rlabel metal2 s 22176 0 22232 400 6 wbs_dat_i[5]
port 337 nsew signal input
rlabel metal2 s 24864 0 24920 400 6 wbs_dat_i[6]
port 338 nsew signal input
rlabel metal2 s 27552 0 27608 400 6 wbs_dat_i[7]
port 339 nsew signal input
rlabel metal2 s 30240 0 30296 400 6 wbs_dat_i[8]
port 340 nsew signal input
rlabel metal2 s 32928 0 32984 400 6 wbs_dat_i[9]
port 341 nsew signal input
rlabel metal2 s 9632 0 9688 400 6 wbs_dat_o[0]
port 342 nsew signal output
rlabel metal2 s 36512 0 36568 400 6 wbs_dat_o[10]
port 343 nsew signal output
rlabel metal2 s 39200 0 39256 400 6 wbs_dat_o[11]
port 344 nsew signal output
rlabel metal2 s 41888 0 41944 400 6 wbs_dat_o[12]
port 345 nsew signal output
rlabel metal2 s 44576 0 44632 400 6 wbs_dat_o[13]
port 346 nsew signal output
rlabel metal2 s 47264 0 47320 400 6 wbs_dat_o[14]
port 347 nsew signal output
rlabel metal2 s 49952 0 50008 400 6 wbs_dat_o[15]
port 348 nsew signal output
rlabel metal2 s 52640 0 52696 400 6 wbs_dat_o[16]
port 349 nsew signal output
rlabel metal2 s 55328 0 55384 400 6 wbs_dat_o[17]
port 350 nsew signal output
rlabel metal2 s 58016 0 58072 400 6 wbs_dat_o[18]
port 351 nsew signal output
rlabel metal2 s 60704 0 60760 400 6 wbs_dat_o[19]
port 352 nsew signal output
rlabel metal2 s 12320 0 12376 400 6 wbs_dat_o[1]
port 353 nsew signal output
rlabel metal2 s 63392 0 63448 400 6 wbs_dat_o[20]
port 354 nsew signal output
rlabel metal2 s 66080 0 66136 400 6 wbs_dat_o[21]
port 355 nsew signal output
rlabel metal2 s 68768 0 68824 400 6 wbs_dat_o[22]
port 356 nsew signal output
rlabel metal2 s 71456 0 71512 400 6 wbs_dat_o[23]
port 357 nsew signal output
rlabel metal2 s 74144 0 74200 400 6 wbs_dat_o[24]
port 358 nsew signal output
rlabel metal2 s 76832 0 76888 400 6 wbs_dat_o[25]
port 359 nsew signal output
rlabel metal2 s 79520 0 79576 400 6 wbs_dat_o[26]
port 360 nsew signal output
rlabel metal2 s 82208 0 82264 400 6 wbs_dat_o[27]
port 361 nsew signal output
rlabel metal2 s 84896 0 84952 400 6 wbs_dat_o[28]
port 362 nsew signal output
rlabel metal2 s 87584 0 87640 400 6 wbs_dat_o[29]
port 363 nsew signal output
rlabel metal2 s 15008 0 15064 400 6 wbs_dat_o[2]
port 364 nsew signal output
rlabel metal2 s 90272 0 90328 400 6 wbs_dat_o[30]
port 365 nsew signal output
rlabel metal2 s 92960 0 93016 400 6 wbs_dat_o[31]
port 366 nsew signal output
rlabel metal2 s 17696 0 17752 400 6 wbs_dat_o[3]
port 367 nsew signal output
rlabel metal2 s 20384 0 20440 400 6 wbs_dat_o[4]
port 368 nsew signal output
rlabel metal2 s 23072 0 23128 400 6 wbs_dat_o[5]
port 369 nsew signal output
rlabel metal2 s 25760 0 25816 400 6 wbs_dat_o[6]
port 370 nsew signal output
rlabel metal2 s 28448 0 28504 400 6 wbs_dat_o[7]
port 371 nsew signal output
rlabel metal2 s 31136 0 31192 400 6 wbs_dat_o[8]
port 372 nsew signal output
rlabel metal2 s 33824 0 33880 400 6 wbs_dat_o[9]
port 373 nsew signal output
rlabel metal2 s 6048 0 6104 400 6 wbs_stb_i
port 374 nsew signal input
rlabel metal2 s 6944 0 7000 400 6 wbs_we_i
port 375 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 110000 75000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 15100446
string GDS_FILE /run/media/tholin/d9eb5833-69bc-462f-98fb-b7c5c019399b/AS2650/openlane/wrapped_as2650/runs/23_11_23_15_26/results/signoff/wrapped_as2650.magic.gds
string GDS_START 532814
<< end >>

