* NGSPICE file created from wrapped_as2650.ext - technology: gf180mcuC

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_2 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_4 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_64 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_64 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_32 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_32 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fill_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fill_1 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_4 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__antenna abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__antenna I VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xnor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xnor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_16 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__fillcap_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__fillcap_8 VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_1 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__filltie abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__filltie VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_16 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_1 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_1 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux2_2 I0 I1 S Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_1 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_1 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_1 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkinv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkinv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi21_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi21_2 A1 A2 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_1 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_3 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__endcap abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__endcap VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_4 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or2_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or2_1 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_2 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai31_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai31_1 A1 A2 A3 B ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_4 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nand2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nand2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor4_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor4_2 A1 A2 A3 A4 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_2 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi221_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi221_1 A1 A2 B1 B2 C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__inv_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__inv_1 I ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__or3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__or3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__clkbuf_8 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_2 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_2 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and4_1 A1 A2 A3 A4 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__and3_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__and3_1 A1 A2 A3 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor3_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor3_4 A1 A2 A3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_2 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tiel abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tiel ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__buf_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__buf_2 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_2 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__tieh abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__tieh Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyc_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyc_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi222_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi222_1 A1 A2 B1 B2 C1 C2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dlyb_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dlyb_1 I Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__mux4_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__mux4_1 I0 I1 I2 I3 S0 S1 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__nor2_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__nor2_4 A1 A2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__dffq_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__dffq_2 D CLK Q VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi211_4 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi211_4 A1 A2 B C ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__xor2_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__xor2_2 A1 A2 Z VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__aoi22_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__aoi22_2 A1 A2 B1 B2 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai33_1 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai33_1 A1 A2 A3 B1 B2 B3 ZN VDD VSS
.ends

* Black-box entry subcircuit for gf180mcu_fd_sc_mcu7t5v0__oai32_2 abstract view
.subckt gf180mcu_fd_sc_mcu7t5v0__oai32_2 A1 A2 A3 B1 B2 ZN VDD VSS
.ends

.subckt wrapped_as2650 io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ vdd vss wb_clk_i wb_rst_i
XFILLER_67_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6914_ _2659_ _2877_ _2890_ _2747_ _2891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_23_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6845_ _2796_ _2822_ _2823_ _2824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_4
XFILLER_126_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6776_ _2046_ _2699_ _2044_ _2047_ _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5196__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3988_ _3501_ _3522_ _3523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_108_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5727_ _0662_ _1746_ _1755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4943__A2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6160__I _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6145__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5658_ _3433_ _1695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4609_ _0758_ _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5589_ _3556_ _1628_ _0422_ _1629_ _1630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_117_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7328_ _0139_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7259_ _0070_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5120__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output37_I net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3959__I _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A2 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4934__A2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3737__A3 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6136__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6136__B2 _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7404__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5111__A2 _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_60_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_64_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4960_ _3209_ _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3911_ as2650.addr_buff\[5\] _3387_ _3446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_60_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4891_ _0929_ _1005_ _1006_ _0937_ _1007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_71_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6630_ _1508_ _1510_ _2615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3842_ _3345_ _3355_ _3376_ _3377_ _3378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_34_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6561_ as2650.psl\[5\] _2459_ _2561_ _2562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4925__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3773_ _3308_ _3241_ _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5512_ _1554_ _1547_ _1556_ _0158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6492_ _2490_ _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5443_ _3142_ _1495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5374_ _1433_ _1434_ _1435_ _1436_ _1437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__5350__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7113_ _0445_ _0974_ _3058_ _3064_ _3065_ _3066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4325_ _0446_ _0521_ _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7044_ _3009_ _2989_ _3011_ _0235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_101_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4256_ as2650.holding_reg\[5\] _3246_ _0454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5102__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4187_ _0374_ _0385_ _0386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6602__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A3 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4613__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6828_ _2680_ _2791_ _2807_ _2640_ _2808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5927__C _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6366__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6759_ _3566_ _3570_ _3541_ _2741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_17_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7427__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5234__I _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__B1 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6774__B _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4852__A1 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_73_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4604__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A2 _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5837__C _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6109__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6949__B _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4110_ _3164_ _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7085__A2 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5090_ _3256_ _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4983__I _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6832__A2 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4041_ _3299_ _3460_ _3489_ _3575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_110_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3646__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5992_ _1324_ _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4943_ _1046_ _1053_ _1056_ _1057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6348__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4874_ _0483_ _0883_ _0990_ _0991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_18_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6613_ _0717_ _2602_ _2605_ _0210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3825_ _3359_ _3360_ _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6544_ _2541_ _0394_ _2542_ _2545_ _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_140_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3756_ as2650.r123\[1\]\[0\] as2650.r123_2\[1\]\[0\] as2650.psl\[4\] _3292_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_14_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6475_ _1506_ _1342_ _2480_ _2481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3687_ _3204_ _3205_ _3212_ _3222_ _3223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_106_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5426_ _1482_ _0146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6520__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5357_ _1419_ _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4308_ _0361_ _0505_ _0506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5288_ _1374_ _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6594__B _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__B1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7027_ _2997_ _3529_ _2998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4239_ _3494_ _0437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6823__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5229__I _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4133__I _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5562__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3876__A2 _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7067__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5899__I _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4825__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6578__A1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6578__B2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4053__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5567__C _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3610_ _3144_ _3145_ _3146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6750__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4590_ as2650.stack\[3\]\[1\] _0761_ _0763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4978__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__B _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3882__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6260_ _2043_ _2096_ _2098_ _2270_ _2271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_127_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6502__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5211_ _1317_ _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_43_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6191_ as2650.stack\[5\]\[6\] _1975_ _2079_ as2650.stack\[4\]\[6\] _2204_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5856__A3 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5142_ as2650.psl\[7\] _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_123_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5073_ _3431_ _3524_ _0274_ _0961_ _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4024_ _3543_ _3467_ _3468_ _3557_ _3558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_49_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__B1 _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4218__I _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6569__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7272__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5975_ as2650.pc\[1\] _3462_ _1992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_0_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4926_ _1031_ _1039_ _1040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4857_ as2650.r0\[4\] _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3808_ _3168_ _3278_ _3344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5544__A2 _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6741__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4788_ _0866_ _0910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6589__B _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6741__B2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6527_ _1685_ _0325_ _2530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3739_ _3180_ _3146_ _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6458_ _1225_ _2463_ _2464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5409_ as2650.stack_ptr\[1\] _1457_ _1470_ _1471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6389_ _1781_ _2395_ _2396_ _1639_ _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__7049__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6608__I _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6009__B1 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6771__C _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5232__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4035__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6980__A1 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__A2 _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3794__A1 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6799__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5422__I _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7295__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4274__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4026__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5760_ _1786_ _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4711_ _0813_ _0838_ _0843_ _0070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5691_ _0368_ _1723_ _1701_ _1724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_7430_ _0241_ clknet_leaf_0_wb_clk_i as2650.r123\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4642_ as2650.stack\[2\]\[7\] _0792_ _0796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6723__A1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5526__A2 _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7361_ _0172_ clknet_leaf_6_wb_clk_i as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4573_ _0747_ _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6312_ _2321_ _1453_ _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7292_ _0103_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6243_ _2254_ _2255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6856__C _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6174_ _2154_ _2155_ _2186_ _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_48_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A3 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5125_ _3466_ _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5332__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5056_ _0668_ _0884_ _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_55_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4007_ _3540_ _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6591__C _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3787__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5214__A1 _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6163__I _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5958_ _1971_ _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5765__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3776__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4909_ _0597_ _0921_ _1024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5889_ _1154_ _1753_ _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5517__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__C _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6714__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6190__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5242__I _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_10_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__A1 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4256__A2 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_57_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6953__A1 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A2 _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_14_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_138_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6181__A2 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5417__I _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4192__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4192__B2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5861__B _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6248__I _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5152__I _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5039__A4 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5444__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6930_ net35 _2905_ _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_66_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6861_ _1776_ _2182_ _2645_ _2839_ _2840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5812_ _1779_ _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6792_ _2770_ _2771_ _2772_ _2773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6944__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5743_ _1586_ _1760_ _1770_ _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_124_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5674_ _1696_ _1697_ _1699_ _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_30_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7413_ _0224_ clknet_leaf_28_wb_clk_i net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4625_ _0783_ _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7344_ _0155_ clknet_leaf_13_wb_clk_i as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4183__A1 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4556_ _0733_ _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7275_ _0086_ clknet_leaf_62_wb_clk_i as2650.r123_2\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_1_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7121__A1 _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4487_ _0669_ _0673_ _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6226_ _2009_ _2226_ _2237_ _3222_ _2238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_89_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6475__A3 _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4387__B _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5683__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6157_ _2132_ _2140_ _2170_ _2037_ _2171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5108_ _1218_ _0989_ _1221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6088_ _1989_ _2102_ _1997_ _2103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5286__I1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4238__A2 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5039_ _3175_ _3357_ _1150_ _1151_ _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XTAP_2705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3997__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5738__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6935__A1 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6935__B2 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4410__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6621__I _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5237__I _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4141__I _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xoutput20 net20 io_out[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_122_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7112__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput31 net31 io_out[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput42 net42 io_out[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6466__A3 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4229__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7179__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7333__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6926__B2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5575__C _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5147__I _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4165__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4410_ _0551_ _0543_ _0605_ _0606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5390_ _1452_ _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5901__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3912__A1 _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4341_ _0396_ _0372_ _0459_ _0496_ _0538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4986__I _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7103__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7060_ _3023_ _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4272_ _0263_ _3552_ _0283_ _0340_ _0470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_87_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6011_ as2650.stack\[7\]\[2\] _1968_ _2027_ as2650.stack\[4\]\[2\] _2028_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_113_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6090__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6913_ _2449_ _2883_ _2889_ _2628_ _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_54_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4226__I _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6844_ _1099_ _0474_ _2823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_126_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6775_ _2625_ _2755_ _2756_ _0221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3987_ _3422_ _3503_ _3519_ _3521_ _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XANTENNA__6393__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6441__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5726_ _1258_ _1753_ _1754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5657_ _1488_ _1692_ _1693_ _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_4608_ _0759_ _0773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5588_ _3171_ _3173_ _3370_ _3476_ _1629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_102_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3903__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4539_ as2650.pc\[6\] _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7327_ _0138_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7258_ _0069_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7206__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5656__A1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6209_ _0720_ _0715_ _2131_ _2221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7189_ _0000_ clknet_leaf_2_wb_clk_i as2650.r123\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_58_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7356__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4136__I _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4631__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4395__A1 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3737__A4 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6136__A2 _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4147__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4622__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3910_ _3353_ _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4890_ _0547_ _0935_ _1006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3841_ _3317_ _3377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4386__A1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6560_ _1049_ _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3772_ _3303_ _3305_ _3307_ _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_5511_ _1555_ _1549_ _1556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_73_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6491_ _1115_ _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5442_ _1054_ _1493_ _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7229__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5373_ _0672_ _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7112_ _0308_ _0961_ _3065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4324_ _0455_ _0520_ _0521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5638__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7043_ _0975_ _2991_ _2992_ _3010_ _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_99_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4255_ _3506_ _0446_ _0451_ _0452_ _0453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7379__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4186_ _3580_ _0384_ _0289_ _0286_ _0385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_83_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4861__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5810__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3996__S _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_23_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6827_ _2638_ _2793_ _2806_ _1831_ _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3795__I _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6171__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6758_ _1298_ _0331_ _2740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_137_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5709_ _1736_ _1737_ _1738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_104_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6689_ _3465_ _3449_ _2672_ _2673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__5943__C _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5877__A1 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5629__A1 _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5629__B2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5250__I _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6054__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__A2 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3654__B _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5868__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6293__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4040_ _3299_ _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_49_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5160__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6045__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5991_ _2007_ _1988_ _1055_ _2008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6596__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4942_ _1055_ _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6348__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4873_ _0480_ _0886_ _0888_ _0990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6205__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4504__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6612_ as2650.stack\[7\]\[5\] _2603_ _2605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3824_ _3180_ _3148_ _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3755_ as2650.r123\[0\]\[0\] as2650.r123_2\[0\]\[0\] as2650.psl\[4\] _3291_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_6543_ _2541_ _2543_ _2544_ _2545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3686_ _3221_ _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6474_ _3174_ _3316_ _3262_ _2480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5859__A1 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5425_ as2650.r123_2\[0\]\[3\] _0972_ _1480_ _1482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4531__A1 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5356_ _3266_ _0656_ _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4307_ _0504_ _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5287_ _1377_ _0112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5087__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__I1 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4238_ _0367_ _0434_ _0436_ _0004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7026_ _2990_ _2997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4395__B _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4169_ as2650.holding_reg\[4\] _0368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5070__I _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5003__C _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4598__A1 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4414__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5245__I _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_39_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6275__A1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A1 as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6578__A2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5848__C _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6750__A2 net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5583__C _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5210_ _3274_ _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_48_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4513__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6190_ as2650.stack\[7\]\[6\] _2164_ _1977_ as2650.stack\[6\]\[6\] _2203_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_142_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5141_ _1117_ _1182_ _1253_ _1116_ _0090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4994__I _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6266__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5072_ _1183_ _1184_ _1185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_38_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4023_ _3469_ _3556_ _3557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6018__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6018__B2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7417__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4943__B _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6569__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5974_ _0699_ _1239_ _1991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4925_ _1034_ _1038_ _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_127_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4856_ _0393_ _0974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3807_ _3342_ _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_140_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6741__A2 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4787_ _0907_ _0908_ _0909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4752__A1 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6526_ _2517_ _0331_ _2529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3738_ _3148_ _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6457_ _2458_ _3343_ _2460_ _2462_ _2463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_133_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3669_ _3195_ _3200_ _3205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5408_ _1469_ _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6388_ _1781_ _2377_ _2396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5339_ as2650.stack\[5\]\[7\] _1404_ _1408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6257__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7009_ net38 _2654_ _1461_ _2982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4853__B _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5232__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output12_I net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6980__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4144__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4743__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5299__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6496__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5703__I _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6799__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6420__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6971__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4710_ as2650.stack\[0\]\[2\] _0839_ _0843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A1 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5690_ _1721_ _1722_ _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4989__I _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6184__B1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4641_ _0722_ _0791_ _0795_ _0048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4572_ as2650.pc\[12\] _0747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7360_ _0171_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6311_ as2650.addr_buff\[1\] _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7291_ _0102_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6487__A1 _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6487__B2 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6242_ as2650.stack\[3\]\[7\] _0649_ _1924_ as2650.stack\[2\]\[7\] _2254_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6173_ _1099_ _0407_ _2186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5613__I _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5124_ _0879_ _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5055_ _0869_ _0358_ _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6872__C _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4006_ _3539_ _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5769__B _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6444__I _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4392__C _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5214__A2 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_52_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5957_ _1970_ _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4908_ _0623_ _0873_ _1020_ _1022_ _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4973__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5888_ _0645_ _1338_ _1907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4839_ _0926_ _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_101_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6509_ _0438_ _3582_ _2513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5009__B _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5523__I _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5453__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6650__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_6_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5205__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6402__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6953__A2 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6166__B1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4016__I0 _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_54_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_4_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7262__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5141__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_45_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6692__C _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5444__A2 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6860_ _1349_ _1418_ _2838_ _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5811_ _1554_ _1153_ _1776_ _1454_ _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_34_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6791_ _2763_ _0330_ _2711_ _2741_ _2742_ _2772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_5742_ _1578_ _1284_ _1765_ _1769_ _1591_ _1770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_124_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5673_ _1708_ _0167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7412_ _0223_ clknet_leaf_28_wb_clk_i net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_124_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4624_ _0784_ _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5904__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7343_ _0154_ clknet_leaf_13_wb_clk_i as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5380__A1 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4555_ as2650.pc\[9\] _0733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_102_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7274_ _0085_ clknet_leaf_0_wb_clk_i as2650.r123_2\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4486_ _0672_ _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7044__B _3011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6439__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6225_ _1652_ _2222_ _2237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_48_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5343__I _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5683__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6156_ _2139_ _2160_ _2169_ _2170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3694__A1 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5107_ _3283_ _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6087_ _2095_ _2094_ _2100_ _2101_ _1995_ _2102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_57_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5038_ _3202_ _1096_ _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_72_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3997__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6989_ _2959_ _2962_ _2963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_15_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__B1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5518__I _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6699__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4422__I _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4174__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xoutput21 net21 io_out[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput32 net32 io_out[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__7112__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput43 net43 io_out[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_123_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6871__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3685__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6623__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3988__A2 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5362__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4165__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4340_ _0536_ _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5114__A1 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4271_ _0468_ _0449_ _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6862__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6010_ _1971_ _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6862__B2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input3_I io_in[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6912_ _1537_ _2888_ _2889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_36_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3979__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6843_ _1099_ _0474_ _2822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_35_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6774_ net28 _2654_ _2694_ _2756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_51_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3986_ _3422_ _3520_ _3521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_22_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5725_ _1752_ _1631_ _1753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3600__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5656_ _3311_ _1259_ _1693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4607_ _0772_ _0037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5587_ _3536_ _0348_ _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7326_ _0137_ clknet_leaf_37_wb_clk_i as2650.stack\[5\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__A2 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4538_ _0718_ _0712_ _0719_ _0021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7257_ _0068_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4469_ _3215_ _0655_ _3213_ _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5656__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6853__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6208_ _1799_ _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7188_ _3128_ _3130_ _2496_ _0260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_86_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6139_ _1269_ _2110_ _2153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6605__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6081__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4092__A1 _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7097__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4101__B _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5647__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6844__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5711__I _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3840_ _3366_ _3370_ _3371_ _3375_ _3376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4386__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5583__A1 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5158__I _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3771_ _3306_ _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4062__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5510_ _0659_ _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6490_ _2493_ _2495_ _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_34_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5441_ _0660_ _1492_ _1493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4138__A2 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5335__A1 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5372_ _1054_ _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7111_ _3059_ _3062_ _3063_ _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7088__A1 _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4323_ _3259_ _0417_ _0519_ _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5638__A2 _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7042_ _2993_ _0500_ _3010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4254_ _0375_ _0377_ _0389_ _0440_ _0450_ _0452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_99_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4310__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4185_ _0284_ _0384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4074__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7012__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6452__I _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6826_ _2799_ _2805_ _1677_ _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_144_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4377__A2 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5574__A1 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6757_ _2665_ _2737_ _2738_ _2667_ _2739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3969_ _3418_ _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5708_ _1729_ _1155_ _3237_ _1737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6688_ _3372_ _3390_ _2672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_137_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5326__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4129__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5639_ _1618_ _1677_ _1678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4700__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5877__A2 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3888__A1 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7079__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7309_ _0120_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7323__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5629__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5531__I _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output42_I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6054__A2 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A1 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5801__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3812__A1 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4368__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5565__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5868__A2 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3879__A1 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6817__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6045__A2 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5990_ _1337_ _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4056__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4941_ _1054_ _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3896__I _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4872_ _0497_ _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6611_ _0710_ _2602_ _2604_ _0209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3823_ _3144_ _3145_ _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5556__A1 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6542_ _2452_ _0400_ _2544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3754_ _3289_ _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_53_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_9_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_9_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__3845__B _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6473_ _1052_ _1065_ _1086_ _1121_ _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_3685_ _3214_ _3220_ _3221_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4520__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5424_ _1481_ _0145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5355_ _1417_ _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4531__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4306_ _3389_ _0418_ _0469_ _0327_ _0503_ _0504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5286_ as2650.r123_2\[1\]\[1\] _0942_ _1375_ _1377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_59_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6284__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7025_ _2990_ _2996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4237_ as2650.r123\[2\]\[4\] _0435_ _0436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4295__A1 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4168_ _3289_ _0367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4099_ _3582_ _3588_ _0288_ _0298_ _0299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_15_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A1 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6809_ _2097_ _2758_ _2789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6744__B1 _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5970__B _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6275__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5261__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4286__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6027__A2 net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4806__S _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7219__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4589__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__A1 net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4210__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6976__B _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4513__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6695__C _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5140_ _1202_ _1252_ _1182_ _1253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_97_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6266__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5069__A3 _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_29_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5071_ _0596_ _1184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4022_ _3546_ _3555_ _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_96_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6018__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5777__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5973_ _1940_ _1990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6216__B _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4515__I _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4924_ _3137_ _1037_ _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5529__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4855_ _0973_ _0084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3806_ _3319_ _3340_ _3341_ _3342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4786_ _0872_ _0908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6525_ _2527_ _2528_ _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7047__B _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3737_ _3253_ _3256_ _3239_ _3272_ _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_107_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6456_ as2650.carry _2461_ _2458_ _2462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3668_ _3203_ _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5407_ _1459_ _1469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5701__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6387_ _2392_ _2394_ _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3599_ _3134_ _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5338_ _0823_ _1403_ _1407_ _0133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6257__A2 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4268__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5269_ _0850_ _1361_ _1366_ _0105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7008_ _2976_ _2980_ _2981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_75_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_68_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6009__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5768__A1 _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A1 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6640__I _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4743__A2 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6796__B _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6496__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4259__A1 _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4806__I0 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6420__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7191__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4982__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4640_ as2650.stack\[2\]\[6\] _0792_ _0795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6184__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6184__B2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4571_ _0745_ _0736_ _0746_ _0027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5931__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6310_ _2009_ _2306_ _2233_ _2320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7290_ _0101_ clknet_leaf_44_wb_clk_i as2650.stack\[6\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6241_ _1971_ _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6172_ _2176_ _2183_ _2184_ _2185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5115__B _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6239__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5123_ _0559_ _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5054_ _3204_ _1166_ _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5998__A1 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4005_ _3538_ _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_72_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5956_ as2650.stack\[3\]\[1\] _1968_ _1969_ as2650.stack\[2\]\[1\] _1973_ _1974_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4907_ _0908_ _1021_ _1022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_142_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5887_ _1149_ _1905_ _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4973__A2 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6175__A1 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4838_ _0274_ _0867_ _0957_ _0958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_14_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5922__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4769_ _0879_ _0883_ _0890_ _0891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_88_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6508_ _2496_ _2498_ _2512_ _0198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_101_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__C _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6439_ _1744_ _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5289__I0 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5989__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_4_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4155__I _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3994__I as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4964__A2 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6370__I _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6166__A1 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4016__I1 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4716__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5913__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7407__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7134__C _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5141__A2 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5444__A3 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4652__A1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5810_ _1832_ _1833_ _1834_ _0657_ _1835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6790_ _1270_ _0406_ _2771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4404__A1 _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5741_ _1105_ _0687_ _1767_ _1768_ _1769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_96_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5672_ _3502_ _1707_ _1701_ _1708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6157__A1 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6157__B2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7411_ _0222_ clknet_leaf_27_wb_clk_i net29 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4623_ _0783_ _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7342_ _0153_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4554_ _0732_ _0024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5380__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7273_ _0084_ clknet_leaf_64_wb_clk_i as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5624__I _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4485_ _0671_ _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6224_ _2233_ _2234_ _2235_ _2236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_131_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5132__A2 _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6155_ _1743_ _2132_ _2168_ _1919_ _2169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3694__A2 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5106_ _1097_ _1209_ _1217_ _1218_ _1219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6086_ _1914_ _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6093__B1 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6455__I _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6632__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5037_ _3254_ _1049_ _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_100_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4643__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_14_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6396__A1 as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6988_ _2413_ _2837_ _2961_ _2870_ _1939_ _2962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_0_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5939_ net2 _1956_ _1957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_139_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4703__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6148__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6148__B2 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_31_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5962__C _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput11 net11 io_oeb[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5534__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xoutput22 net22 io_out[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput33 net33 io_out[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput44 net44 io_out[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3685__A2 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4882__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6365__I _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6623__A2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6387__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4937__A2 _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6139__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5898__B1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5362__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4270_ _0395_ _0370_ _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5114__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6984__B _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6862__A2 _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3676__A2 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6614__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6911_ _2885_ _2887_ _2888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6842_ net32 _2820_ _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6378__A1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6773_ _2041_ _2658_ _2754_ _2692_ _2755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_62_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3985_ _3502_ _3355_ _3419_ _3520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5050__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5724_ _1603_ _1752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3600__A2 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5655_ _1266_ _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_opt_4_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6878__C _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4606_ _0731_ as2650.stack\[3\]\[8\] _0759_ _0772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5586_ _1602_ _1605_ _1626_ _1627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_7325_ _0136_ clknet_leaf_35_wb_clk_i as2650.stack\[5\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4537_ as2650.stack\[4\]\[5\] _0713_ _0719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5354__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6302__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7256_ _0067_ clknet_leaf_38_wb_clk_i as2650.stack\[1\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4468_ _3216_ _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_131_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6207_ as2650.pc\[7\] _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7187_ _1694_ _3108_ _3129_ _3130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_113_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4399_ _3398_ _0594_ _0595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4864__A1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6138_ _1269_ _2110_ _2152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6605__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6069_ as2650.stack\[2\]\[3\] _2078_ _2084_ as2650.stack\[0\]\[3\] _2085_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_3227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3602__I _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4616__A1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__B1 _1836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_139_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5592__A2 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4147__A3 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7097__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6844__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4608__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3770_ as2650.idx_ctrl\[1\] as2650.idx_ctrl\[0\] _3306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5583__A2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5440_ _0661_ _0684_ _1492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6532__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5371_ _0668_ _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7110_ _0274_ _3061_ _3063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4322_ _0447_ _0262_ _0519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7088__A2 _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7041_ net41 _3009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6835__A2 _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4253_ _0375_ _0377_ _0450_ _0451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_68_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4846__A1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4184_ _3512_ _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7275__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4074__A2 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_3_7_0_wb_clk_i clknet_0_wb_clk_i clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__7012__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6825_ _2674_ _2803_ _2804_ _2715_ _2805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5023__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6771__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3968_ _3502_ _3354_ _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5574__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6756_ _0345_ _2476_ _2738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6889__B _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6771__B2 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5793__B _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5707_ _1460_ _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6687_ _2670_ _2671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3899_ _3432_ _3433_ _3434_ _3272_ _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_136_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5638_ _1675_ _1676_ _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6523__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5326__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5569_ _1558_ _1152_ _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3888__A2 _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7308_ _0119_ clknet_leaf_56_wb_clk_i as2650.r123\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7079__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7239_ _0050_ clknet_leaf_39_wb_clk_i as2650.stack\[2\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5812__I _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4837__A1 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output35_I net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4065__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5262__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6643__I _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_42_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_14_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5565__A2 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6514__A1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3879__A2 _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6817__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7298__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6039__B _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4056__A2 _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6553__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4940_ _3147_ _3219_ _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4871_ _0988_ _0085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6610_ as2650.stack\[7\]\[4\] _2603_ _2604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3822_ _3356_ _3357_ _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6753__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5556__A2 _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6541_ _2450_ _0406_ _2543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3753_ _3138_ _3288_ _3289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6505__A1 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6472_ _3303_ _0379_ _1168_ _1657_ _2478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
X_3684_ _3215_ _3217_ _3219_ _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_88_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5423_ as2650.r123_2\[0\]\[2\] _0958_ _1480_ _1481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_106_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5354_ _1416_ _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4305_ _0328_ _0471_ _0503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5285_ _1376_ _0111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7024_ _2983_ _2989_ _2995_ _0231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4236_ _3439_ _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4167_ _3290_ _0365_ _0366_ _0003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5788__B _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4098_ _0270_ _0265_ _0298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__A1 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5795__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6992__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6808_ _2657_ _2788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6744__A1 _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6744__B2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6739_ _2004_ _2698_ _2005_ _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5807__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7440__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6638__I _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4038__A2 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6432__B1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A1 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_48_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4822__S _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6735__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5717__I _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4210__A2 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4621__I _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3721__A1 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5070_ _3264_ _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_78_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5474__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4068__I _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4021_ _3547_ _3548_ _3472_ _3554_ _3555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__3901__S _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4029__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5777__A2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3700__I _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5972_ _1889_ _1989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6216__C _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4923_ _1035_ _1036_ _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_94_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5529__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4854_ _0972_ as2650.r123_2\[2\]\[3\] _0959_ _0973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_60_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3805_ as2650.psl\[3\] as2650.carry _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4785_ _3391_ _0878_ _0906_ _0907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6524_ _1710_ _2494_ _1736_ _2528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3736_ _3265_ _3271_ _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7151__A1 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6455_ _1873_ _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3667_ _3202_ _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5406_ _1464_ _1467_ _1468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6386_ _0686_ _2278_ _2393_ _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3598_ as2650.ins_reg\[0\] _3134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5337_ as2650.stack\[5\]\[6\] _1404_ _1407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5268_ as2650.stack\[6\]\[7\] _1362_ _1366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_9_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6662__B1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7007_ _0748_ _2657_ _2979_ _1939_ _2726_ _2980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_4219_ _0417_ _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5199_ _1306_ _1309_ _1310_ _1311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5217__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__A2 _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3779__A1 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4440__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5965__C _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3703__A1 _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5272__I _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5205__C _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5456__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7336__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6956__A1 net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4431__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6184__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4570_ as2650.stack\[4\]\[11\] _0737_ _0746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5931__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7133__A1 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6240_ _1970_ _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6171_ _1799_ _2184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5122_ _0483_ _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_97_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5447__A1 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5053_ _3207_ _3356_ _3211_ _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_69_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5998__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5910__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4004_ net3 _3538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_65_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6947__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5955_ _1972_ _1973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4906_ _0603_ _0947_ _1021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5886_ _1895_ _1901_ _1904_ _1905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_16_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4973__A3 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4837_ _0944_ _0956_ _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5357__I _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6175__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4261__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4768_ _3370_ _0886_ _0889_ _0890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5922__A2 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6507_ _0892_ _1855_ _2502_ _2503_ _2511_ _2512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7124__A1 _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3719_ _3254_ _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5293__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4699_ _0749_ _0828_ _0834_ _0067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6438_ _0748_ _1883_ _2443_ _2444_ _1595_ _0196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__7209__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5092__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6369_ as2650.pc\[11\] _2376_ _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5438__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__C _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4436__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5610__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6166__A2 net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4177__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4171__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4104__C _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7115__A1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_63_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_63_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4346__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4652__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4790__B _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5601__B2 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5740_ _1555_ _1636_ _1763_ _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5671_ _1704_ _1706_ _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5177__I _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4081__I as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7410_ _0221_ clknet_leaf_27_wb_clk_i net28 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4622_ _0757_ _0782_ _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5904__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7341_ _0152_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4553_ _0731_ as2650.stack\[4\]\[8\] _0691_ _0732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_144_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5905__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7272_ _0083_ clknet_leaf_64_wb_clk_i as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4484_ _3138_ _3405_ _0670_ _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_132_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5668__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6223_ _1268_ _1416_ _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4030__B _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6154_ _2163_ _2167_ _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5105_ _1048_ _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6085_ _2097_ _2099_ _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6093__B2 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5036_ _1034_ _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6632__A3 _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5840__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5691__I1 _1723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6987_ _2392_ _2446_ _2960_ _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6396__A2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5938_ as2650.r123\[2\]\[1\] as2650.r123_2\[2\]\[1\] _3324_ _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5869_ _1426_ _1423_ _1775_ _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6148__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4159__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__A1 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput12 net12 io_oeb[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput23 net23 io_out[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput34 net34 io_out[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xoutput45 net45 io_out[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4882__A2 _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6084__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6387__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4398__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3996__I1 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6139__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5898__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5898__B2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5362__A3 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5114__A3 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7161__B _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3676__A3 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4873__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__A1 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6075__B2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_82_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6910_ _3307_ _2886_ _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_35_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6841_ net51 _2792_ _2820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6378__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4389__A1 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6772_ _2542_ _2750_ _2753_ _2050_ _2754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3984_ _3511_ _3518_ _3519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5050__A2 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5723_ _1489_ _0685_ _1424_ _1665_ _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5654_ _3185_ _1687_ _1690_ _1691_ _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5889__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4605_ _0726_ _0766_ _0771_ _0036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6550__A2 _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5585_ _1611_ _1625_ _1626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4561__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7324_ _0135_ clknet_leaf_44_wb_clk_i as2650.stack\[5\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4536_ _0717_ _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7255_ _0066_ clknet_leaf_37_wb_clk_i as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4467_ _3206_ _3361_ _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_131_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6206_ _0722_ _1936_ _2218_ _0190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4398_ _3423_ _0575_ _0594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7186_ _3114_ _1693_ _3129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4864__A2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6137_ _1512_ _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5370__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6068_ _0804_ _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4616__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5813__B2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5019_ _1123_ _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4714__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_127_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5545__I _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4147__A4 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6541__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7097__A3 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4304__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_27_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6057__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A1 _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_opt_4_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_83_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6325__B _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4624__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4791__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4543__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5370_ _1324_ _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4321_ _0514_ _0517_ _0518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7088__A3 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6296__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7040_ _3002_ _3007_ _3008_ _0234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4252_ _0447_ _0449_ _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_87_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_141_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4183_ _0300_ _0378_ _0381_ _3408_ _0382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_67_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7012__A3 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6824_ _1101_ _2674_ _2804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6220__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6755_ _0344_ _0325_ _2736_ _2737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3967_ as2650.holding_reg\[1\] _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6771__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5706_ _0576_ _1727_ _1735_ _0173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4782__A1 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6686_ _2669_ _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3898_ _3239_ _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_34_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5637_ _3224_ _1495_ _1497_ _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6523__A2 _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5731__B1 _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5568_ _1048_ _1177_ _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7307_ _0118_ clknet_leaf_62_wb_clk_i as2650.r123_2\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4519_ _0702_ _0692_ _0703_ _0018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5499_ _1535_ _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3814__S _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6287__A1 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7238_ _0049_ clknet_leaf_36_wb_clk_i as2650.stack\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4837__A2 _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7169_ _3113_ _3115_ _3116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_98_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6039__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5262__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6145__B _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6211__A1 as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4773__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6514__A2 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6278__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__B2 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6450__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5253__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_75_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4870_ _0987_ as2650.r123_2\[2\]\[4\] _0959_ _0988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3821_ _3156_ _3210_ _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_53_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6540_ _1201_ _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4764__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3752_ _3287_ _3288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6502__C _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6471_ _3184_ _2476_ _1129_ _2477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3683_ _3218_ as2650.cycle\[0\] _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5185__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5422_ _1476_ _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_86_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5353_ _3270_ _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4304_ _0476_ _3484_ _0499_ _0501_ _3315_ _0502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_114_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5284_ as2650.r123_2\[1\]\[0\] _0912_ _1375_ _1376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7242__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4529__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7023_ _3311_ _2991_ _2992_ _2994_ _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4235_ _3496_ _0394_ _0433_ _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_25_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4166_ as2650.r123\[2\]\[3\] _3440_ _0366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4097_ _0294_ _0295_ _0296_ _0297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_83_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5244__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5795__A3 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__I1 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6807_ _2625_ _2785_ _2787_ _0222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6744__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4999_ _1096_ _1112_ _1113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6738_ _1056_ _1344_ _2720_ _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_136_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6669_ _2623_ _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5483__A2 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6680__A1 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6654__I _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6432__A1 as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3797__A2 _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6735__A2 _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_17_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_17_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6499__A1 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7265__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5171__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3721__A2 _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4349__I _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6671__A1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4020_ _3549_ _3553_ _3554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5474__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6423__A1 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4029__A3 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5971_ _1986_ _1987_ _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4922_ as2650.psl\[7\] _0676_ _1036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4853_ _0961_ _0867_ _0971_ _0972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6726__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3804_ _3339_ _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4784_ _0891_ _0898_ _0905_ _0906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_18_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6523_ _2497_ _2520_ _2525_ _2526_ _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_140_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3735_ _3270_ _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3960__A2 _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6454_ as2650.psu\[0\] _2459_ _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3666_ _3153_ _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_133_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__A1 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5405_ _1466_ _0651_ _0755_ _1467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6385_ as2650.addr_buff\[0\] _2321_ as2650.addr_buff\[2\] _2393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
X_3597_ _3132_ _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5336_ _0821_ _1403_ _1406_ _0132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5267_ _0823_ _1361_ _1365_ _0104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_29_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6662__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7006_ as2650.pc\[12\] _2684_ _2978_ _2870_ _2432_ _2979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5799__B _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6662__B2 _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4218_ _0416_ _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5198_ _1033_ _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4149_ _0346_ _0348_ _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5217__A2 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6965__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5768__A3 _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3779__A2 _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4722__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7288__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_109_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7142__A2 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5153__A1 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6350__B1 _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4900__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5456__A2 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6384__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6405__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_74_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4719__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3942__A2 _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7133__A2 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5144__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6170_ _2095_ _2175_ _2182_ _2101_ _1995_ _2183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_139_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5121_ _0425_ _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5052_ _0356_ _3168_ _1165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_85_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6294__I as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4003_ _3536_ _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3711__I _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4958__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5954_ as2650.stack\[1\]\[1\] _1970_ _1971_ as2650.stack\[0\]\[1\] _1972_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_0_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4905_ _0948_ _1018_ _1019_ _0947_ _1020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__7430__CLK clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5885_ _1893_ _1902_ _1903_ _1509_ _1904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_80_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__A1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4836_ _3577_ _0946_ _0955_ _0956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5383__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4767_ _0888_ _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6506_ _2491_ _2510_ _2511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3718_ _3158_ _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7124__A2 _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4698_ as2650.stack\[1\]\[12\] _0829_ _0834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5135__A1 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6437_ _1885_ _2415_ _1935_ _2444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_135_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5373__I _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3649_ as2650.idx_ctrl\[1\] _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_103_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6368_ _0739_ _2340_ _2376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5319_ _0689_ _0806_ _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6299_ _0728_ _1280_ _2309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5438__A2 _1419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6635__A1 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5610__A2 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5374__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4177__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7115__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5283__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6874__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7303__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6328__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7051__A1 net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5601__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4362__I _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_32_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5670_ _3483_ _1705_ _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6998__B _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4621_ _0781_ _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5365__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7340_ _0151_ clknet_leaf_14_wb_clk_i as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_11_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4552_ _0730_ _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7106__A2 _3522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6314__B1 _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7271_ _0082_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4483_ _3202_ _3178_ _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6865__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6222_ _0659_ _1806_ _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5668__A2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_49_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6153_ _2030_ _2165_ _2166_ _2167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_112_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5921__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5104_ _0868_ _1210_ _1108_ _1216_ _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_98_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6084_ _2043_ _2098_ _2099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_111_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5035_ _0358_ _1141_ _1147_ _1053_ _1148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_73_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5840__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__C _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6986_ _2445_ _2953_ _2960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5937_ net1 _3293_ _1955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5368__I _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3603__A1 as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5868_ _0646_ _1885_ _1886_ _1887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5356__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4819_ _0908_ _0939_ _0940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4159__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5799_ _0655_ _3219_ _3268_ _1824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3906__A2 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6420__C _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5108__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3616__I _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7326__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput13 net13 io_oeb[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5659__A2 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xoutput24 net24 io_out[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
Xoutput35 net35 io_out[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_27_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_102_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6084__A2 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XPHY_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6847__A1 _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5114__A4 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6837__I _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6058__B _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5897__B _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6840_ _2178_ _2818_ _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_78_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5035__B1 _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6771_ _2041_ _2684_ _2752_ _1428_ _1257_ _2753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_126_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4389__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5586__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3983_ _3512_ _3514_ _3515_ _3516_ _3517_ _3518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_108_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5722_ _1039_ _1749_ _1746_ _1750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_50_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5338__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5653_ _1575_ _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6535__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7349__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4604_ as2650.stack\[3\]\[7\] _0767_ _0771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4010__A1 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5584_ _1614_ _1615_ _1616_ _1624_ _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_7_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7323_ _0134_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4535_ _0716_ _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4041__B _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7254_ _0065_ clknet_leaf_37_wb_clk_i as2650.stack\[1\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4466_ _3140_ _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_132_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3880__B _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6205_ _2130_ _2216_ _2217_ _2218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4313__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5651__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7185_ as2650.psu\[0\] _3127_ _3128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4397_ _0588_ _0591_ _0592_ _3423_ _0593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6136_ _2066_ _2145_ _2148_ _2149_ _2150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6067_ as2650.stack\[3\]\[3\] _2075_ _2082_ as2650.stack\[1\]\[3\] _2083_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4077__A1 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5018_ _1060_ _1107_ _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3824__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7015__A1 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5577__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6969_ _2933_ _2939_ _2943_ _1205_ _2944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_42_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5329__A1 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4001__A1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6829__A1 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5804__A2 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3815__A1 as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7006__B2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5568__A1 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5736__I _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4791__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4543__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5672__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4320_ _0515_ _0516_ _0517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7088__A4 _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7172__B _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4288__S _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4251_ _0448_ _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5471__I _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4182_ _0379_ _0341_ _0380_ _0300_ _0381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA_input1_I io_in[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__B _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_51_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5559__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6823_ _0482_ _0505_ _2802_ _2803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_90_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4606__I0 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5023__A3 _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6754_ _2704_ _2734_ _2735_ _2736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3966_ _3397_ _3500_ _3501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4231__A1 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5705_ _1727_ _1734_ _1735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6685_ as2650.addr_buff\[7\] _3230_ _2669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__4782__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3897_ _3303_ _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5646__I _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5636_ _1528_ _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_12_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6523__A3 _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5567_ _1258_ _1066_ _1516_ _1564_ _1607_ _1608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5731__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5731__B2 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7306_ _0117_ clknet_leaf_62_wb_clk_i as2650.r123_2\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4518_ as2650.stack\[4\]\[2\] _0693_ _0703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_2_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5498_ _1544_ _1536_ _1546_ _0154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6287__A2 _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7237_ _0048_ clknet_leaf_39_wb_clk_i as2650.stack\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4449_ as2650.r123\[1\]\[5\] _0637_ _0639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5381__I _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7168_ _3114_ _1721_ _1722_ _3115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6039__A2 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6119_ as2650.pc\[5\] net6 _2133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7099_ _1741_ _0394_ _3039_ _3040_ _3052_ _3053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_74_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5798__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4725__I _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A1 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5970__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4773__A2 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4460__I _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5722__A1 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6278__A2 _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4289__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3804__I _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4635__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6450__A2 _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4461__A1 as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6055__C _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3820_ _3163_ _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4213__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3751_ _3235_ _3252_ _3273_ _3286_ _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_144_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5466__I _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6470_ _3306_ _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3682_ as2650.cycle\[1\] _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5421_ _1479_ _0144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5352_ _0860_ _1410_ _1415_ _0139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6269__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4303_ _3479_ _0500_ _3379_ _0501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5283_ _1374_ _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7022_ _2993_ _3548_ _2994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4234_ _3436_ _0401_ _0432_ _0433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4165_ _3496_ _0315_ _0364_ _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_56_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4096_ _0270_ _0265_ _0285_ _0296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_67_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4452__A1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6806_ net29 _2786_ _2694_ _2787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4998_ _1098_ _1111_ _1112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6737_ _1434_ _0357_ _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3949_ _3312_ _3484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_17_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5376__I _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6668_ _1634_ _2651_ _2652_ _1897_ _2653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_136_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5619_ _1082_ _1321_ _3269_ _0682_ _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_104_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5704__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6599_ _2594_ _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3624__I _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6680__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__C _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_73_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4455__I as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6432__A2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__A1 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5943__B2 _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6499__A2 _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5171__A2 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_57_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_57_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5474__A3 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4682__A1 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6423__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5970_ _0696_ _0644_ _0699_ _1987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4921_ as2650.psl\[6\] _0677_ _1035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6187__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4852_ _0325_ _0873_ _0970_ _0910_ _0971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_100_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3803_ _3338_ _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_127_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5934__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4783_ as2650.r0\[0\] _0900_ _0903_ _3342_ _0904_ _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_92_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5934__B2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6522_ _3556_ _1779_ _1854_ _0332_ _2526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3734_ _3266_ _3181_ _3269_ _3270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_119_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6453_ _1091_ _2459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3665_ _3195_ _3200_ _3201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_118_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5404_ _1465_ _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6384_ as2650.addr_buff\[3\] _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5162__A2 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3596_ _3131_ _3132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_115_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5335_ as2650.stack\[5\]\[5\] _1404_ _1406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5266_ as2650.stack\[6\]\[6\] _1362_ _1365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6111__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7005_ _2428_ _2977_ _2978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6662__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4217_ _0408_ _0409_ _0412_ _0415_ _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_130_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5197_ _1255_ _1307_ _1308_ _1309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_55_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4148_ _3545_ _3554_ _0347_ _0348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_55_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4079_ _0278_ _3396_ _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4425__A1 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5834__I _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6350__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5153__A2 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5456__A3 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_47_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4416__A1 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5916__A1 _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7382__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7164__C _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5144__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_39_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5120_ _1231_ _1232_ _1233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_97_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5051_ _1161_ _1126_ _1163_ _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_112_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4655__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4002_ _3535_ _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_22_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5953_ _0804_ _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5919__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6524__B _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4904_ _0617_ _0948_ _1019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5884_ _3374_ _0664_ _1903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_94_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3630__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4835_ _3571_ _0947_ _0946_ _0954_ _0955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5907__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5907__B2 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6580__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4766_ _0887_ _0888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5383__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6505_ _1834_ _2504_ _2509_ _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3717_ _3195_ _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4697_ _0745_ _0828_ _0833_ _0066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3648_ _3143_ _3182_ _3183_ _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XANTENNA__6332__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6436_ _2434_ _2442_ _1801_ _2443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6367_ _0744_ _2374_ _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__A1 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3697__A2 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5318_ _1394_ _0126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_62_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6298_ _2307_ _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_114_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6485__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6635__A2 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5249_ _1353_ _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_5_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3902__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_2_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5694__I0 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7255__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__A2 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__I1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5374__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6874__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4885__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__B1 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6626__A2 _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4637__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3860__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7159__C _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6011__B1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4620_ _0780_ _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6562__A1 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5365__A2 _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4551_ _0729_ _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7270_ _0081_ clknet_leaf_2_wb_clk_i as2650.r123_2\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5117__A2 _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4482_ _0668_ _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6314__B2 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6221_ _1126_ _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6865__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4876__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6152_ as2650.stack\[2\]\[5\] _1969_ _1975_ as2650.stack\[1\]\[5\] _2166_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5103_ as2650.psl\[6\] _1214_ _1215_ _1216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6617__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6083_ _2046_ _1993_ _2044_ _2047_ _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3722__I _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4628__A1 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5034_ _1142_ _1144_ _1031_ _1146_ _1147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__7278__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4039__B _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7042__A2 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6985_ _1963_ _2385_ _2959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5053__A1 _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5936_ _1157_ _1941_ _1954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3603__A2 net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4800__A1 _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5867_ _1881_ _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5356__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4818_ _3449_ _0878_ _0938_ _0939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4159__A3 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5798_ _3215_ _3217_ _3360_ _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_124_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4749_ _0870_ _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5108__A2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput14 net14 io_oeb[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput25 net25 io_out[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6856__A2 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6419_ _1898_ _2415_ _2426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xoutput36 net36 io_out[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7399_ _0210_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__B1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4728__I _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3632__I _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3842__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7033__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4463__I _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7420__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5035__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5035__B2 _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_0 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6770_ _1418_ _2733_ _2751_ _2752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3982_ _3404_ _3164_ _3517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5586__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5721_ _1163_ _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3918__S _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__A1 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5652_ _3229_ _1689_ _1687_ _1690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6535__B2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4603_ _0722_ _0766_ _0770_ _0035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5583_ _1617_ _1619_ _1620_ _1623_ _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_117_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3717__I _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4534_ _0715_ _0716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_116_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7322_ _0133_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_85_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7253_ _0064_ clknet_leaf_38_wb_clk_i as2650.stack\[1\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4465_ as2650.stack_ptr\[2\] _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6204_ _1469_ _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7184_ _1237_ _1733_ _3108_ _3127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4396_ _0576_ _3420_ _3340_ _0592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6135_ _1102_ _1513_ _1815_ _3228_ _1258_ _2149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6066_ _0780_ _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5017_ _0676_ _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_38_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4283__I net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6968_ _2373_ _2684_ _2942_ _2644_ _2943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_53_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5919_ as2650.pc\[1\] _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6899_ _2858_ _2859_ _2876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5329__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3627__I _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7443__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5265__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3815__A2 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7006__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5568__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_38_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6517__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5238__B _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3981__B _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5752__I _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4250_ _0408_ _0409_ _0412_ _0415_ _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_114_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4181_ _0368_ _0379_ _0380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3806__A2 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4854__I1 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5008__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7316__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6822_ _2770_ _2800_ _2772_ _2801_ _2802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XANTENNA__5559__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6756__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6753_ _3540_ _3573_ _3576_ _2735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_32_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3965_ _3499_ _3500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4231__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5704_ _1554_ _1733_ _1267_ _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6508__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3896_ _3253_ _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6684_ _2662_ _2664_ _2666_ _2667_ _2668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_31_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3990__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__B _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5635_ _1662_ _1673_ _1674_ _1576_ _0163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_136_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5566_ _1083_ _1524_ _1341_ _1606_ _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XANTENNA__5731__A2 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7305_ _0116_ clknet_leaf_62_wb_clk_i as2650.r123_2\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3742__A1 _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4517_ _0701_ _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5497_ _1545_ _1538_ _1546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7236_ _0047_ clknet_leaf_40_wb_clk_i as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4448_ _0434_ _0636_ _0638_ _0012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4278__I as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4379_ as2650.holding_reg\[7\] _0574_ _0575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7167_ _1109_ _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6118_ _0716_ _2131_ _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7098_ _3050_ _3051_ _3052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5247__A1 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_86_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6049_ _1525_ _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3910__I _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6995__A1 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6426__C _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4470__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4222__A2 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4741__I _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3981__A1 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5722__A2 _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__A1 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5572__I _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4289__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5238__A1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4916__I _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7339__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6986__A1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4461__A2 as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5747__I _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3750_ _3278_ _3285_ _3286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4764__A3 _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5961__A2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3681_ _3216_ _3217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__7163__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7163__B2 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5420_ as2650.r123_2\[0\]\[1\] _0942_ _1477_ _1479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_9_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6910__A1 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5351_ as2650.stack\[5\]\[12\] _1411_ _1415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4302_ _0342_ _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5282_ _1061_ _0925_ _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4233_ _3384_ _0406_ _0431_ _3442_ _0432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7021_ _2990_ _2993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4164_ _3436_ _0326_ _0363_ _0364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_68_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4826__I _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3730__I _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4095_ _3581_ _0287_ _0295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_67_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_fanout52_I net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6729__A1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6805_ _2623_ _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_24_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4997_ as2650.psu\[5\] _1103_ _1105_ _1110_ _1111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_6736_ _1501_ _2698_ _2700_ _1786_ _2718_ _2719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3948_ _3482_ _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_71_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6667_ _1850_ _1689_ _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7154__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3879_ _3395_ _3406_ _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5165__B1 _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5618_ _0863_ _1160_ _1168_ _1657_ _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6901__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5704__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6598_ _2595_ _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6488__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7093__B _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3715__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5392__I _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5549_ _1203_ _1518_ _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_2_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__A1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7219_ _0030_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4140__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5483__A4 _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3640__I _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__B2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4443__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_54_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5943__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3954__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7145__A1 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3706__A1 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_29_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_6_0_wb_clk_i clknet_0_wb_clk_i clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_124_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__B1 _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_0_wb_clk_i_I wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5474__A4 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4682__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4646__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5631__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_52_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4920_ _1033_ _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4851_ _0872_ _0969_ _0970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_2690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6187__A2 _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4198__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3802_ _3337_ _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4782_ _3382_ _0871_ _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6521_ _1229_ _2523_ _2524_ _2525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3733_ _3268_ _3217_ _3213_ _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__7136__A1 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6452_ _1218_ _2458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3664_ _3199_ _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5403_ _1439_ _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6383_ _1802_ _2379_ _2390_ _2391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3595_ as2650.ins_reg\[1\] _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5162__A3 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4370__A1 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5334_ _0817_ _1403_ _1405_ _0131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5265_ _0821_ _1361_ _1364_ _0103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6111__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7004_ _1745_ _2967_ _2977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4122__A1 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4216_ _0333_ as2650.r123\[1\]\[5\] _3326_ _0414_ _0415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5196_ _1042_ _1045_ _1308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4147_ _3281_ _3368_ _3354_ _3545_ _0347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_95_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4078_ _3395_ _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5622__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4425__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4189__A1 _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_7_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6719_ _3462_ _3491_ _2702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5689__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6350__A2 _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3635__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6102__A2 _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4113__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4664__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5861__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4466__I _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6681__I _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5916__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7118__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7017__I _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5760__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4104__A1 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5050_ _1027_ _1106_ _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4001_ _3532_ _3534_ _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5852__A1 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A1 net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5952_ _0780_ _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_18_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4903_ _0989_ _0918_ _1017_ _0895_ _1018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_80_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5883_ _1488_ _3293_ _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_61_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3630__A3 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4834_ _0948_ _0952_ _0953_ _0937_ _0954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_14_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4765_ _3175_ _3167_ _0874_ _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__7109__B2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6504_ _1292_ _1232_ _2507_ _2508_ _1587_ _2509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_135_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4591__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3716_ _3236_ _3241_ _3251_ _3252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_88_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4696_ as2650.stack\[1\]\[11\] _0829_ _0833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6435_ _1918_ _2416_ _2441_ _2442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3647_ as2650.cycle\[6\] _3145_ _3183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_134_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6366_ _2373_ _2352_ _2374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4894__A2 _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5317_ as2650.r123\[3\]\[7\] _1394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6297_ _0733_ _1211_ _2307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_142_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6096__A1 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5248_ _0689_ _0782_ _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6635__A3 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5694__I1 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5843__A1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5179_ _3373_ _1291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_56_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4949__A3 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6450__B _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5374__A3 _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6571__A2 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4582__A1 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4885__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__B2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5062__A2 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6011__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__B _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4550_ _0728_ _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4481_ _3279_ _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5691__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6220_ _0725_ _2231_ _2232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_144_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5704__B _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4876__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_41_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_41_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6151_ as2650.stack\[3\]\[5\] _2164_ _1976_ as2650.stack\[0\]\[5\] _2165_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6078__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__C _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5102_ _1173_ _1214_ _1215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6082_ _2096_ _2097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4628__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5033_ _1145_ _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6984_ _2861_ _2957_ _2866_ _2958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_25_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6250__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__A2 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5935_ _1775_ _1938_ _1943_ _1908_ _1952_ _1953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5866_ _1884_ _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6002__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4817_ _0929_ _0934_ _0936_ _0937_ _0938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_33_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5797_ _1797_ _0655_ _1798_ _1822_ _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4748_ _3253_ _0869_ _3139_ _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_108_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6305__A2 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4679_ as2650.stack\[1\]\[5\] _0819_ _0822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4316__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6418_ _2423_ _2424_ _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
Xoutput15 net15 io_oeb[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput26 net52 io_out[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_7398_ _0209_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput37 net37 io_out[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6349_ _1890_ _2356_ _2357_ _2358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_89_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7222__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5816__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4619__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_48_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7372__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6544__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_45_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6480__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6232__A1 net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5035__A2 _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_1 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_1_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3981_ _3502_ _3248_ _3405_ _3516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_62_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6783__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5720_ _1745_ _1635_ _1746_ _1747_ _1748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_50_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4794__A1 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__C _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5651_ _1613_ _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5485__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6535__A2 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4602_ as2650.stack\[3\]\[6\] _0767_ _0770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5582_ _1584_ _1622_ _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7321_ _0132_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4533_ as2650.pc\[5\] _0715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7252_ _0063_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4464_ _0650_ _0651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7245__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6203_ _2175_ _2185_ _2214_ _2215_ _2216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7183_ _3124_ _3126_ _0259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_131_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4395_ _3408_ _0590_ _0444_ _0591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6249__C _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6134_ _1056_ _2146_ _2147_ _2148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5153__C _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7395__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6065_ _2024_ _2077_ _2080_ _2081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_100_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6471__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5016_ _1125_ _1128_ _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4564__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7015__A3 _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6223__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5026__A2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6967_ _1344_ _2346_ _2645_ _2941_ _2942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_53_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6774__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4785__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5918_ _1935_ _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6898_ _2816_ _2873_ _2875_ _0225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5849_ _1607_ _1864_ _1867_ _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5395__I _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3908__I _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6526__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4537__A1 as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_120_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_67_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6462__A1 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4474__I _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4776__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3818__I _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7268__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7025__I _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4180_ _3248_ _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5256__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6205__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6821_ _0423_ _0405_ _2801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6756__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6752_ _3573_ _3576_ _3540_ _2734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3964_ _3258_ _3471_ _3498_ _3499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5703_ _1259_ _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6683_ _2627_ _2667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3895_ _3430_ _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4519__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5634_ net22 _1662_ _1674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3990__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7181__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5192__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5565_ _1047_ _1080_ _1081_ _1606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7304_ _0115_ clknet_leaf_3_wb_clk_i as2650.r123_2\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4516_ _0700_ _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3742__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5496_ as2650.addr_buff\[3\] _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7235_ _0046_ clknet_leaf_40_wb_clk_i as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4559__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4447_ as2650.r123\[1\]\[4\] _0637_ _0638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7166_ _3088_ _3112_ _3113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_86_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4378_ _3320_ _3322_ _3330_ _3336_ _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_98_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6117_ _0709_ _0704_ _1986_ _2131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XTAP_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7097_ _1103_ _1692_ _1150_ _3051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5247__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6048_ _1811_ _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5798__A3 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6995__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6723__B _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4758__A1 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7410__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3638__I _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3981__A2 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7172__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_19_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5722__A3 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4930__A1 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5238__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6435__A1 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_40_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6986__A2 _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__B _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6738__A2 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4764__A4 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3811__I3 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3972__A2 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3680_ as2650.cycle\[2\] _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7163__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5174__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6371__B1 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5350_ _0858_ _1410_ _1414_ _0138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4301_ _0485_ _0498_ _0499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5281_ _0860_ _1368_ _1373_ _0110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7020_ _2988_ _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4232_ _0429_ _0430_ _0361_ _0431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_64_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4163_ _3384_ _0331_ _0362_ _3442_ _0363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_95_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6426__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6426__B2 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4094_ _3591_ _3509_ _0293_ _0294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_95_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7433__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6729__A2 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6804_ _2135_ _2652_ _2784_ _1634_ _2785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_24_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4996_ _1102_ _1109_ _1110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6735_ _2701_ _2717_ _2718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3947_ as2650.r0\[1\] _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6666_ _2642_ _2650_ _2651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3963__A2 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3878_ _3413_ _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5165__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5617_ _3316_ _1155_ _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5165__B2 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6597_ _2594_ _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6901__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5548_ _1587_ _1589_ _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_3_0_wb_clk_i clknet_3_6_0_wb_clk_i clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_105_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5479_ _0864_ _1530_ _1531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6665__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5468__A2 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7218_ _0029_ clknet_leaf_24_wb_clk_i as2650.stack\[3\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_99_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7149_ _3319_ _3098_ _3099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4140__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__A1 as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6968__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7090__A1 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4979__A1 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5640__A2 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output26_I net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout50 net34 net50 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_23_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6353__B1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4903__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4903__B2 _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7306__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6656__A1 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__B2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_2_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3831__I _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7081__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6423__A4 _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5631__A2 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6363__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4662__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4850_ _0331_ _0878_ _0968_ _0969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3801_ _3320_ _3322_ _3330_ _3336_ _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4198__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4781_ _0902_ _0899_ _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5694__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6520_ _3543_ _1229_ _1078_ _2524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3732_ _3267_ _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3945__A2 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6451_ _1263_ _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3663_ _3197_ _3198_ _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5402_ _0651_ _0755_ _1463_ _1464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6382_ _1566_ _1424_ _2387_ _2389_ _2390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_103_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3594_ net23 net18 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_86_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5162__A4 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5333_ as2650.stack\[5\]\[4\] _1404_ _1405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4370__A2 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5264_ as2650.stack\[6\]\[5\] _1362_ _1364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7003_ _2971_ _2975_ _2976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_87_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4215_ _3192_ _0413_ _0414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5195_ _0611_ _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_60_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4146_ _0317_ _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__B _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7072__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4077_ _3290_ _0276_ _0277_ _0002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4572__I as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5386__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4189__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4979_ _1050_ _1090_ _1092_ _1093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_138_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6718_ _1676_ _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5138__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6649_ _3391_ _2633_ _2634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3916__I _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7329__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5689__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4113__A2 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5861__A2 _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6810__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5578__I _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4482__I _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A1 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7118__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3826__I _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6877__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6341__A3 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6358__B _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5301__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4104__A2 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4000_ _3198_ _3533_ _3534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5604__A2 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6801__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5951_ _0753_ _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4902_ _0613_ _0915_ _1016_ _1017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5882_ _1431_ _1900_ _1901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4833_ _3528_ _0935_ _0953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_107_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6565__B1 _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4764_ _3169_ _0884_ _0885_ _0870_ _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_140_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6503_ _3283_ _3451_ _0332_ _1088_ _1263_ _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3715_ _3244_ _3250_ _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_105_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4591__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4695_ _0831_ _0828_ _0832_ _0065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6434_ _1919_ _2437_ _2440_ _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3646_ _3180_ _3181_ _3182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_140_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6365_ _2339_ _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5316_ _1393_ _0125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_66_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6296_ _2304_ _2305_ _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_27_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6096__A2 _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5247_ _3356_ _1331_ _1352_ _0097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_9_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5178_ net24 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__3854__A1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6782__I _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4129_ _0328_ _0321_ _0322_ _0329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_56_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5398__I _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4949__A4 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5374__A4 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4582__A2 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6859__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4477__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6087__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__B _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3845__A1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5810__B _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4270__A1 _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3757__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6011__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4022__A1 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5770__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4480_ _3256_ _0278_ _3242_ _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_144_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5771__I _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6150_ _1967_ _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6078__A2 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5101_ _1213_ _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_32_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6081_ _0708_ net5 _2096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5032_ _3362_ _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_leaf_10_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_10_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6535__C _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5589__A1 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6983_ _2380_ _2956_ _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6250__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5053__A3 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6107__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5934_ _1944_ _1945_ _1951_ _1430_ _1952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_20_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5011__I _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5865_ _0864_ _1613_ _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6551__B _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6002__A2 _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4816_ _0876_ _0937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4013__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5796_ _1801_ _1820_ _1821_ _1619_ _1774_ _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_119_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5761__A1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4071__B _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4747_ _0336_ _0868_ _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_108_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4678_ _0717_ _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6417_ as2650.pc\[12\] _1280_ _2424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_134_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5513__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3629_ _3160_ _3164_ _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7397_ _0208_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5681__I _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput16 net16 io_oeb[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput27 net27 io_out[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_1_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput38 net38 io_out[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6348_ _1433_ _2341_ _2357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6069__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6279_ _2054_ _2281_ _2289_ _1424_ _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5816__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3827__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6687__I _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__A1 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7009__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7197__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4491__A1 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6232__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3980_ _3260_ _3355_ _3515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5291__I0 as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_62_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5991__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4794__A2 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4670__I _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5650_ _3186_ _1687_ _1688_ _1576_ _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_15_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4601_ _0718_ _0766_ _0769_ _0034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5743__A1 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5581_ _1621_ _1139_ _1154_ _1622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7320_ _0131_ clknet_leaf_42_wb_clk_i as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_106_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4532_ _0711_ _0712_ _0714_ _0020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_8_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6299__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7251_ _0062_ clknet_leaf_40_wb_clk_i as2650.stack\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6597__I _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4463_ _0649_ _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6202_ _1800_ _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7182_ as2650.psu\[1\] _3125_ _1461_ _3126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4394_ _0578_ _0589_ _0590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6133_ _1653_ _2132_ _2147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6064_ as2650.stack\[6\]\[3\] _2078_ _2079_ as2650.stack\[4\]\[3\] _2080_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5015_ _1126_ _1127_ _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6471__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6223__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5026__A3 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6966_ _1542_ _2191_ _2940_ _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4234__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5917_ _1882_ _1935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6897_ net33 _2786_ _2874_ _2875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_21_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5848_ _1517_ _1579_ _1866_ _1032_ _1663_ _1867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_139_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5734__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4537__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5779_ _1802_ _1665_ _1804_ _1805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7449_ _0260_ clknet_leaf_7_wb_clk_i as2650.psu\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3924__I _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4755__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6462__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_72_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_48_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4776__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4490__I _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3751__A3 _3273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_99_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_113_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7041__I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6820_ _0423_ _0405_ _2800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4216__A1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6751_ net28 _2732_ _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3963_ _3497_ _3257_ _3498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5964__A1 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5496__I as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5702_ _1727_ _1731_ _1732_ _0172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6682_ _1238_ _2665_ _2666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3894_ _3398_ _3402_ _3426_ _3429_ _3430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_91_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7212__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5633_ _1663_ _1672_ _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4519__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5564_ _1175_ _1604_ _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5192__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4515_ _0699_ _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7303_ _0114_ clknet_leaf_64_wb_clk_i as2650.r123_2\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5495_ _1298_ _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7362__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6141__A1 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4446_ _0630_ _0637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7234_ _0045_ clknet_leaf_46_wb_clk_i as2650.stack\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7165_ _3107_ _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4377_ _0367_ _0572_ _0573_ _0006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6116_ _1882_ _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7096_ _3046_ _3049_ _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6047_ _2056_ _2062_ _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4758__A2 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6949_ _1537_ _1540_ _2482_ _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4016__S _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6380__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_5_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3733__A3 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4930__A2 _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4485__I _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4997__A2 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_4_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6633__C _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7235__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5946__A1 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__C1 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7385__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__A1 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__A2 _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6371__B2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4921__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4300_ _3345_ _0497_ _3377_ _0498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6123__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5280_ as2650.stack\[6\]\[12\] _1369_ _1373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4231_ as2650.r0\[4\] _0359_ _0430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4685__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4162_ _0353_ _0360_ _0361_ _0362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_96_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6426__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4093_ _3499_ _3583_ _0293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6803_ _2455_ _2778_ _2783_ _2784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5937__A1 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4995_ _0869_ _1108_ _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6734_ _2708_ _2716_ _2717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3946_ _3450_ _3451_ _3480_ _3481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6665_ _1785_ _2649_ _2650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3877_ _3399_ _3401_ _3413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5616_ _1623_ _1648_ _1650_ _1655_ _1656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6362__A1 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6362__B2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6596_ _0689_ _0755_ _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5547_ _1588_ _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6114__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5478_ _1529_ _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_144_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6665__A2 _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4429_ _3443_ _0620_ _0624_ _3494_ _0625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7217_ _0028_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4676__A1 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7148_ _3092_ _3097_ _3098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6417__A2 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7079_ _0653_ _1319_ _3035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7258__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7090__A2 _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4979__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3651__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A1 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6025__I as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout51 net31 net51 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4600__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5864__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6353__B2 as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_89_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6105__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6656__A2 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3800_ _3194_ as2650.r123\[0\]\[7\] _3333_ _3335_ _3336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
X_4780_ _0901_ _3282_ _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3731_ as2650.cycle\[3\] _3267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_119_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_35_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5774__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6344__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3662_ as2650.ins_reg\[0\] _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6450_ _2056_ _3431_ _2455_ _2456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5401_ _1142_ _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6381_ as2650.addr_buff\[3\] _1512_ _2388_ _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_103_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5332_ _1395_ _1404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5723__B _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6647__A2 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5263_ _0817_ _1361_ _1363_ _0102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7002_ _1832_ _2973_ _2974_ _2975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4214_ as2650.r123_2\[1\]\[5\] _0413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_114_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5194_ _1046_ _1304_ _1305_ _1306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_96_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4145_ _0344_ _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5014__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3881__A2 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4076_ as2650.r123\[2\]\[2\] _3440_ _0277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6554__B _2217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5083__A1 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5949__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4830__A1 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5386__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6583__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4978_ _1091_ _1092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6717_ _1991_ _2699_ _2700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_20_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3929_ _3463_ _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6335__A1 as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5138__A2 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6648_ _2632_ _2633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6579_ _2576_ _2578_ _1232_ _2579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4897__A1 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4649__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7063__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5074__A1 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6810__A2 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4821__A1 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5377__A2 _1038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5594__I _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6326__A1 _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4888__A1 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4003__I _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7423__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6629__A2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5301__A2 _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7054__A2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5065__A1 _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4673__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6801__A2 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5950_ _1967_ _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_94_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6093__C _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4812__A1 _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4901_ _0607_ _0978_ _0915_ _1015_ _1016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_5881_ _1433_ _1896_ _1899_ _1435_ _1900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6014__B1 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4832_ _0892_ _0918_ _0951_ _0952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6565__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6565__B2 _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4763_ _3214_ _3220_ _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_18_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6502_ as2650.psu\[1\] _2505_ _2506_ _1090_ _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6317__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3714_ _3249_ _3250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4694_ as2650.stack\[1\]\[10\] _0829_ _0832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6868__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6433_ _1922_ _2438_ _2439_ _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3645_ as2650.cycle\[0\] _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_128_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4879__A1 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6364_ _0741_ _1936_ _2372_ _0194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5453__B _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5315_ as2650.r123\[3\]\[6\] _1393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7371__D _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6295_ _0728_ _2263_ _2305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3752__I _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5246_ _1351_ _1339_ _1352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5177_ _1270_ _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4128_ _3385_ as2650.addr_buff\[6\] _0328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__A1 _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4059_ _3581_ _3592_ _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_71_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__A1 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A1 _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3927__I net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6308__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7446__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6859__A2 _2821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3790__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3863__S _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3662__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4098__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7036__A2 _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5810__C _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__I0 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6244__B1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6795__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3999__I3 as2650.r123_2\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4270__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6547__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5538__B _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3837__I _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5770__A2 _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3781__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5100_ _1212_ _1213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6080_ _1940_ _2095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XTAP_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4089__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6883__I _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5031_ _1143_ _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7027__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5499__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5038__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6982_ _2381_ _2936_ _2956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5589__A2 _1628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6786__A1 _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5933_ _1133_ _1950_ _1124_ _1951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_0_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_50_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_59_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5864_ _1882_ _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4815_ _3482_ _0935_ _0936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7366__D _0177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5795_ _3251_ _1657_ _1698_ _1808_ _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4746_ _3135_ _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3772__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4677_ _0817_ _0818_ _0820_ _0059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6416_ _2420_ _2421_ _2422_ _2423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5513__A2 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3628_ _3161_ _3163_ _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7396_ _0207_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput17 net17 io_oeb[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_134_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput28 net28 io_out[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_116_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput39 net39 io_out[2] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6347_ _2007_ _2346_ _2356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6278_ _2230_ _2283_ _2288_ _1075_ _2289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_83_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5277__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5229_ _1337_ _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3827__A2 _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_38_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4252__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5201__A1 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3763__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5872__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6701__A1 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5504__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4488__I _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_140_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5268__A1 as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6465__B1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6480__A3 _1151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4491__A2 _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6208__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6768__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5112__I _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5440__A1 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_3 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4951__I _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5991__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4600_ as2650.stack\[3\]\[5\] _0767_ _0769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5743__A2 _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5580_ _3209_ _1118_ _1621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_89_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4531_ as2650.stack\[4\]\[4\] _0713_ _0714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7250_ _0061_ clknet_leaf_40_wb_clk_i as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4462_ _0648_ _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6201_ _2183_ _2200_ _2213_ _2214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4393_ _0515_ _0513_ _0516_ _0532_ _0589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_7181_ _3102_ _3112_ _3125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6132_ _1338_ _2138_ _2146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__B _2806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6063_ _0804_ _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5014_ _0663_ _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6471__A3 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A1 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6965_ _2151_ _2931_ _2940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5957__I _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5916_ _0646_ _1883_ _1887_ _1934_ _1853_ _0184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_35_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6896_ _1459_ _2874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3993__A1 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7184__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5847_ _1059_ _1064_ _1865_ _1866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_22_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5778_ _1664_ _3269_ _1803_ _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5734__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3745__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4729_ _0836_ _0855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4810__B _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7448_ _0259_ clknet_leaf_54_wb_clk_i as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5498__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7379_ _0190_ clknet_leaf_33_wb_clk_i as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4170__A1 _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5670__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5867__I _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4771__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3984__A1 _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7175__A1 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6922__A1 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5725__A2 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5107__I _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4011__I _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4946__I _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5661__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4681__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6750_ net27 net26 net25 _2732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_17_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3962_ as2650.holding_reg\[1\] _3497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5701_ _0531_ _1727_ _1732_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_92_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6681_ _3307_ _2665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3893_ _3165_ _3427_ _3428_ _3429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5632_ _1664_ _1322_ _1345_ _1554_ _1671_ _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__6913__A1 _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6913__B2 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5563_ _1432_ _1603_ _1604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7302_ _0113_ clknet_leaf_64_wb_clk_i as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4514_ as2650.pc\[2\] _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_89_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5494_ _3543_ _1536_ _1543_ _0153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7233_ _0044_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4445_ _0628_ _0636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6141__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5017__I _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7164_ _1290_ _3109_ _3111_ _3108_ _1595_ _0255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4376_ as2650.r123\[2\]\[6\] _0435_ _0573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6429__B1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6115_ _0711_ _1984_ _2129_ _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3760__I _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7095_ _1514_ _2656_ _3047_ _3048_ _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__6276__C _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6046_ _2059_ _2061_ _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5687__I _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6948_ _2885_ _2887_ _2715_ _2482_ _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3966__A1 _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7157__A1 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6879_ _2850_ _2856_ _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6904__A1 _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6380__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6311__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4391__A1 _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6668__B1 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6132__A2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5891__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4766__I _0887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3670__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__A1 _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5946__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7148__A1 _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5159__B1 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4006__I _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5159__C2 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6371__A2 _2375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6221__I _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6123__A2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4230_ _3318_ _3537_ _0428_ _3379_ _0429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5882__A1 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4161_ _3383_ _0361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4092_ _3408_ _0291_ _0292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_95_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5634__A1 net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4437__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7001__B _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6802_ _2135_ _2721_ _2782_ _2720_ _1204_ _2783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_1_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5937__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4994_ _1107_ _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6733_ _1240_ _2632_ _2714_ _2715_ _2716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3945_ _3452_ _3461_ _3478_ _3479_ _3480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_56_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6664_ _2644_ _2647_ _2648_ _0645_ _2649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_137_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3876_ as2650.psl\[3\] _3411_ _3412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5615_ _1144_ _1651_ _1525_ _1654_ _1655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_118_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6595_ _2587_ _2592_ _2593_ _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_118_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5546_ _1451_ _1557_ _1588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5477_ _1528_ _1498_ _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7216_ _0027_ clknet_leaf_33_wb_clk_i as2650.stack\[4\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4428_ _3488_ _0623_ _0624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5873__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4676__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4586__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7147_ _1715_ _1567_ _3097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4359_ _0552_ _0554_ _0555_ _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_87_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7078_ _0626_ _3029_ _3034_ _0246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_58_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5625__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4428__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6029_ _2043_ _2044_ _2045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_74_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_104_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5210__I _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5928__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4254__C _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3939__A1 _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_3_0_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xfanout52 net26 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_35_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6353__A2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5813__C _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6197__B _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4496__I _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__I0 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7202__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5616__A1 _1623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5631__A4 _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7352__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_90 io_out[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_127_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6592__A2 _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3730_ _3218_ _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_92_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3661_ _3196_ _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5400_ _0751_ _1458_ _1462_ _0140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6380_ _1298_ _1562_ _2233_ _2388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5331_ _1396_ _1403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6819__C _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4107__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__C _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5262_ as2650.stack\[6\]\[4\] _1362_ _1363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7001_ _2661_ _2967_ _2866_ _2974_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5855__A1 _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4213_ _0333_ as2650.r123\[0\]\[5\] _3333_ _0411_ _0412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_102_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5193_ _1254_ _0611_ _0678_ _1108_ _1305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_116_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4144_ _0343_ _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_56_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5607__A1 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4075_ _3496_ _3578_ _0275_ _0276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6280__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5083__A2 _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4830__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5030__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6570__B _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4977_ _1060_ _1074_ _1063_ _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6583__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6716_ _2681_ _1947_ _1992_ _2699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3928_ _3462_ _3463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_32_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6647_ _0658_ _3230_ _2632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6335__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3859_ _3160_ _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6578_ _1223_ _2577_ _0549_ _1220_ _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4897__A2 _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5914__B _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5529_ _1572_ _1449_ _1135_ _1573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A1 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7225__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6271__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5074__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_output31_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6023__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6574__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4337__A1 _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5824__B _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5837__A1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3998__C _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_65_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5065__A2 _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4900_ _1014_ _0978_ _1015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5880_ _1897_ _1898_ _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6014__B2 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4831_ _0346_ _0930_ _0917_ _0950_ _0951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6565__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5785__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4576__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4762_ _3358_ _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6501_ _1279_ _1091_ _2506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3713_ _3171_ _3248_ _3249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6317__A2 _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4693_ _0740_ _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6432_ as2650.stack\[2\]\[12\] _1925_ _2253_ as2650.stack\[0\]\[12\] _2439_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3644_ as2650.cycle\[1\] _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_128_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6363_ _2130_ _2371_ _2217_ _2372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5314_ _1392_ _0124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6294_ as2650.pc\[9\] _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_88_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5245_ _1307_ _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5176_ as2650.psu\[4\] _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4127_ _3386_ _0327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_110_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6253__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5056__A2 _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4058_ _3591_ _3513_ _3503_ _3592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA_clkbuf_leaf_28_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6005__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
Xclkbuf_3_5_0_wb_clk_i clknet_0_wb_clk_i clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_73_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6556__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3790__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4774__I _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6547__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_89_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4014__I _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3781__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5554__B _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6483__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5030_ _1123_ _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7060__I _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6235__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5038__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6981_ _2701_ _2950_ _2954_ _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_20_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5589__A3 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6786__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5932_ _1337_ _1941_ _1949_ _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4797__A1 _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5729__B _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5863_ _1881_ _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_55_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4814_ _0900_ _0935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5794_ _1466_ _1813_ _1817_ _1819_ _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_21_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4745_ _0866_ _0867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5761__A3 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3772__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4676_ as2650.stack\[1\]\[4\] _0819_ _0820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6415_ _0743_ _0558_ _2381_ _2344_ _2422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3627_ _3162_ _3163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7395_ _0206_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xoutput18 net49 io_oeb[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_89_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput29 net29 io_out[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
X_6346_ _1780_ _2354_ _1210_ _2355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4721__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6277_ _1780_ _2285_ _2287_ _2288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6474__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5277__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5228_ _1336_ _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3827__A3 _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_56_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5159_ _1268_ _3339_ _0342_ _1270_ _0419_ _1100_ _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_131_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6226__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6777__A2 _2757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6529__A2 _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_122_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3673__I _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6701__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5268__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6465__B2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4009__I _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5440__A2 _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6940__A2 _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4530_ _0690_ _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4461_ as2650.stack_ptr\[1\] as2650.stack_ptr\[0\] _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_6200_ _2201_ _2175_ _2212_ _2213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7180_ _3102_ _3112_ _3123_ _3124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_113_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4392_ _3506_ _0584_ _0587_ _0383_ _0588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_113_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6131_ _2142_ _2144_ _2145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6827__C _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A1 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5259__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6062_ _0753_ _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5013_ _3362_ _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7436__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6759__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_54_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6964_ _2936_ _2938_ _2640_ _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5915_ _1917_ _1933_ _1801_ _1934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6895_ _2863_ _2867_ _2872_ _2873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7377__D _0188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3993__A2 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5846_ _1621_ _1139_ _1865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7184__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5777_ _0655_ _3219_ _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5973__I _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6392__B1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6931__A2 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_5_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3745__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4728_ _0837_ _0854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7447_ _0258_ clknet_leaf_53_wb_clk_i as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4659_ _0757_ _0806_ _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_11_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6695__A1 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7378_ _0189_ clknet_leaf_33_wb_clk_i as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_66_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6329_ _0735_ _1936_ _2338_ _0193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4170__A2 _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_49_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6998__A2 _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5213__I _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5670__A2 _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3668__I _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7175__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3736__A2 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__B1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6438__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5123__I _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5661__A2 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6663__B _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_29_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_63_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4962__I _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5413__A2 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3961_ _3435_ _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5700_ _1728_ _1729_ _1730_ _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3975__A2 _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6680_ _3465_ _3492_ _2663_ _2664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_3892_ _3397_ _3428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7166__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5631_ net22 _1651_ _1669_ _1670_ _1671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_73_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4924__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5562_ _1069_ _1037_ _1440_ _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_7301_ _0112_ clknet_leaf_1_wb_clk_i as2650.r123_2\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4513_ _0697_ _0692_ _0698_ _0017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5493_ _1542_ _1538_ _1543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6677__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7232_ _0043_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4444_ _0365_ _0629_ _0635_ _0011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7163_ _1728_ _1729_ _3110_ _1236_ _3111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__4152__A2 _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4375_ _0437_ _0537_ _0571_ _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_98_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6557__C _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6114_ _1985_ _2128_ _2039_ _2129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_113_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7094_ _2469_ _1165_ _3048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_28_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6045_ _0343_ _2060_ _2061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5033__I _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5652__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3663__A1 _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5968__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4872__I _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6947_ _2879_ _2881_ _1519_ _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_35_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6878_ _2671_ _2854_ _2855_ _2517_ _2856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_22_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5829_ _1654_ _1850_ _1851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4821__B _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5208__I _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4112__I _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6668__B2 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5652__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5340__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5891__A2 _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7093__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5643__A2 _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3654__A1 _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5878__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5159__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5159__B2 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__B1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4906__A1 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6108__B1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5118__I _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7281__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5562__B _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4957__I _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4160_ _0354_ _0359_ _0360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3893__A1 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7084__A1 _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4091_ _0288_ _0290_ _0291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5634__A2 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6831__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_82_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6801_ _2064_ _2100_ _2781_ _2782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_51_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4993_ _3174_ _0880_ _1106_ _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_90_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6732_ _1500_ _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3944_ _3317_ _3479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4070__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7139__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5737__B _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6663_ _1146_ _1811_ _2643_ _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3875_ as2650.carry _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_108_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6898__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5614_ _1653_ _1434_ _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6594_ _0617_ _2555_ _2569_ _2593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_34_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4373__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5545_ _1455_ _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5476_ _1527_ _1528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4427_ _0622_ _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7215_ _0026_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7390__D _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5873__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7146_ _2496_ _3094_ _3096_ _0252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4358_ _3473_ _0553_ _0543_ _0555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_98_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_8_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7077_ as2650.r123\[0\]\[7\] _3030_ _3034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4289_ _3137_ _0486_ _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5625__A2 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6028_ _0704_ _1297_ _2044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_58_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5698__I _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6338__B1 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4364__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5561__A1 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3681__I _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5616__A2 _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6941__B _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_80 io_oeb[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_91 io_out[36] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6041__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4052__A1 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3660_ as2650.ins_reg\[1\] _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_9_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4355__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5552__A1 _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5330_ _0815_ _1397_ _1402_ _0130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5261_ _1353_ _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_48_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7000_ _2424_ _2972_ _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_4212_ _3192_ _0410_ _0411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5855__A2 _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5192_ _3138_ _1045_ _1287_ _1303_ _1304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_9_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_44_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4143_ net4 _0343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__B2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4074_ _3436_ _0274_ _0275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6280__A2 _2290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4976_ _1089_ _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6715_ net27 _2697_ _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3927_ net2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4594__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3766__I _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3858_ _3302_ _3310_ _3393_ _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6646_ _0879_ _2630_ _2631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5543__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3789_ _3324_ _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_6577_ _0574_ _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5528_ _1257_ _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6099__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4597__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5459_ _1342_ _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5846__A2 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_57_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7129_ _0902_ _1177_ _3046_ _3080_ _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_87_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4282__A1 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output24_I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4034__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5782__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5837__A2 _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_2_0_wb_clk_i clknet_3_5_0_wb_clk_i clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_0_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6014__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4830_ _3556_ _0923_ _0914_ _0949_ _0950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4761_ _0882_ _0883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5773__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7058__I _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3712_ _3247_ _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6500_ _1091_ _2505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_14_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4692_ _0827_ _0828_ _0830_ _0064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3643_ _3178_ _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6431_ as2650.stack\[3\]\[12\] _1929_ _2252_ as2650.stack\[1\]\[12\] _2438_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5525__A1 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6362_ _2341_ _2348_ _2370_ _2215_ _2371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_128_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5313_ as2650.r123\[3\]\[5\] _1392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6293_ _1773_ _2303_ _0192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5244_ _3504_ _1331_ _1350_ _0096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3839__A1 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5175_ _1271_ _1276_ _1286_ _1287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6565__C _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4126_ _3310_ _0325_ _0326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6137__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4057_ _3497_ _3445_ _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_84_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5041__I _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4803__A3 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5764__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4959_ _1061_ _1066_ _1072_ _1052_ _1073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_138_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4319__A2 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5516__A1 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6629_ _0860_ _2609_ _2614_ _0217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5216__I _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7342__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6244__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4255__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5755__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__B _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5507__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3781__A3 _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6180__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4494__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4186__B _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5997__S _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6980_ _2659_ _2953_ _1787_ _2954_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5931_ _1336_ _1948_ _1949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5994__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4797__A2 _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5862_ _1660_ _1868_ _1871_ _1880_ _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7215__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4813_ _3451_ _0903_ _0933_ _0934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5793_ _3220_ _1818_ _1463_ _1819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4744_ _0864_ _3272_ _0865_ _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5745__B _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4675_ _0807_ _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3772__A3 _3307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6414_ _2343_ _2380_ _2421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3626_ as2650.ins_reg\[7\] _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7394_ _0205_ clknet_leaf_49_wb_clk_i as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xoutput19 net19 io_out[0] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_127_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6345_ _2003_ _0687_ _2018_ _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5036__I _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6276_ _1898_ _2264_ _2286_ _1145_ _2287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_115_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A2 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5227_ _3157_ _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_103_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5158_ _1269_ _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_116_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6226__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4109_ _0305_ _0308_ _0309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_110_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4237__A1 as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5089_ _1185_ _1187_ _1198_ _1199_ _1201_ _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_84_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5985__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_72_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_112_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_8_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6162__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4712__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3903__B _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6465__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4476__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7238__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5728__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7388__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4400__A1 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5565__B _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6240__I _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4460_ _0646_ _0647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6153__A1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4391_ _3415_ _0585_ _0586_ _0587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6130_ _0717_ _2143_ _2144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6456__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6061_ as2650.stack\[7\]\[3\] _2075_ _2076_ as2650.stack\[5\]\[3\] _2077_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_97_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4467__A1 _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5012_ _1123_ _1124_ _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6963_ _1786_ _2937_ _2938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_81_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5914_ _1897_ _1918_ _1932_ _1933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6894_ _0725_ _2652_ _2871_ _2215_ _2872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5719__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5845_ _1609_ _1610_ _1864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5776_ _1423_ _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6931__A3 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4727_ _0853_ _0076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3774__I _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7393__D _0204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6144__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7446_ _0257_ clknet_leaf_54_wb_clk_i as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4658_ _0805_ _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6695__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3609_ as2650.cycle\[3\] as2650.cycle\[2\] _3145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7377_ _0188_ clknet_leaf_30_wb_clk_i as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4589_ _0647_ _0760_ _0762_ _0029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6328_ _2130_ _2337_ _2217_ _2338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6447__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6259_ _2134_ _2267_ _2270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_67_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3949__I _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4630__A1 as2650.stack\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6383__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6060__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6135__B2 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4697__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5832__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6438__A2 _1883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5404__I _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3859__I _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6610__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3960_ _3443_ _3487_ _3493_ _3494_ _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4183__C _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3891_ as2650.holding_reg\[0\] _3367_ _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_92_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5630_ _1132_ _1491_ _1670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_34_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6374__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3594__I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4924__A2 _1037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5561_ _1140_ _1601_ _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7300_ _0111_ clknet_leaf_63_wb_clk_i as2650.r123_2\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_121_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4512_ as2650.stack\[4\]\[1\] _0693_ _0698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5492_ as2650.addr_buff\[2\] _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6677__A2 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7231_ _0042_ clknet_leaf_24_wb_clk_i as2650.stack\[2\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4443_ as2650.r123\[1\]\[3\] _0631_ _0635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5742__C _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4374_ _3443_ _0565_ _0570_ _3494_ _0571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_7162_ _1105_ _1109_ _3110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7403__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6429__A2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6113_ _2094_ _2103_ _2127_ _2037_ _2128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7093_ _0913_ _0902_ _3319_ _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6044_ as2650.r123\[2\]\[3\] as2650.r123_2\[2\]\[3\] _3325_ _2060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3663__A2 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7388__D _0199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6601__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6946_ _2816_ _2920_ _2921_ _0227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_74_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4612__A1 as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6877_ _1231_ _2671_ _2855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5828_ _1250_ _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5759_ _1530_ _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6117__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5933__B _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7429_ _0240_ clknet_leaf_3_wb_clk_i as2650.r123\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5425__S _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4679__A1 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7093__A2 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4851__A1 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3654__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4603__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5159__A2 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__A1 as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7426__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3893__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7084__A2 _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4090_ _3580_ _0289_ _0290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6831__A2 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4842__A1 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6800_ _2645_ _2780_ _2781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4992_ _3157_ _3279_ _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6731_ _2711_ _2712_ _2713_ _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3943_ _3466_ _3467_ _3468_ _3477_ _3478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6662_ _1344_ _1896_ _2645_ _2646_ _2647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6347__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3874_ _3403_ _3402_ _3409_ _3410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5613_ _1652_ _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6593_ _0607_ _1837_ _1855_ _2577_ _2591_ _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_125_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5544_ _1577_ _1318_ _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_30_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5570__A2 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5475_ as2650.cycle\[6\] _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7214_ _0025_ clknet_leaf_32_wb_clk_i as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4426_ _3339_ _0316_ _0599_ _3574_ _0621_ _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA_clkbuf_leaf_47_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7145_ _1722_ _3093_ _3095_ _3096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_98_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5044__I _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4357_ _3473_ _0553_ _0538_ _3547_ _0554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_101_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7075__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7076_ _0572_ _3029_ _3033_ _0245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4288_ as2650.r123\[2\]\[6\] as2650.r123_2\[2\]\[6\] _0333_ _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_100_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5086__A1 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6027_ as2650.pc\[3\] net4 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_39_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4833__A1 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5389__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6929_ net50 _2876_ _2905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_39_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6338__B2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7449__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5561__A2 _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6759__B _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__C _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6510__A1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7066__A2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5077__A1 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4793__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_70 io_oeb[26] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_81 io_oeb[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_92 io_out[37] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5838__B _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4052__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6513__I _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5129__I _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4033__I _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5552__A2 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4968__I _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5260_ _1354_ _1361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4211_ as2650.r123_2\[0\]\[5\] _0410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_5191_ _1294_ _1300_ _1302_ _1303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_68_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3866__A2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7057__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4142_ _0341_ _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5068__A1 _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6804__A2 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4073_ _0273_ _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4815__A1 _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_leaf_13_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_13_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_92_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4975_ _1088_ _3283_ _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6714_ net52 net25 _2697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3926_ _3460_ _3461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6645_ _2629_ _3302_ _2630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3857_ _3381_ _3392_ _3310_ _3393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_137_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_34_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6740__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6576_ net24 _2459_ _2575_ _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5543__A2 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6740__B2 _2722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3788_ _3323_ _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6579__B _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_3_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5527_ _1561_ _1564_ _1570_ _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__3782__I _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5458_ _1492_ _1509_ _1510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4099__B _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4409_ _3473_ _0470_ _0459_ _0496_ _0605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_132_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5389_ _1451_ _0662_ _1452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_47_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7128_ _3168_ _1711_ _1695_ _3080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7059_ _3287_ _1042_ _3438_ _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5074__A4 _1186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7271__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5231__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3957__I _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6333__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5782__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3793__A1 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6489__B _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5393__B _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4788__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3692__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_112_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6798__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4273__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5470__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4028__I _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3867__I _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4025__A2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4760_ _3279_ _0881_ _0870_ _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6970__A1 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5773__A2 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6970__B2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3784__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3711_ _3246_ _3247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4691_ as2650.stack\[1\]\[9\] _0829_ _0830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6430_ _1473_ _2435_ _2436_ _2437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3642_ _3170_ _3178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5525__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6722__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6399__B _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6361_ _2347_ _2361_ _2369_ _2370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5312_ _1391_ _0123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7007__C _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6292_ _0730_ _1985_ _2302_ _2303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6486__B1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5243_ _1349_ _1339_ _1350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5174_ _1059_ _1283_ _1284_ _1285_ _1286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_111_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__B1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6238__C2 _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7023__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4125_ _0324_ _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5322__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4056_ _3415_ _3589_ _3590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_71_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3777__I _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4958_ _1067_ _1071_ _1072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5764__A2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3909_ _3383_ _3444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5992__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4889_ _0463_ _0918_ _1003_ _1004_ _1005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_119_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6628_ as2650.stack\[7\]\[12\] _2610_ _2614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5516__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6559_ _1466_ _0480_ _2560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_105_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6477__B1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5452__A1 _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5204__A1 _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6952__A1 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5755__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6704__A1 _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5507__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6704__B2 _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6180__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5407__I _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4191__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6947__B _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4494__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4246__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5930_ _1946_ _1947_ _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_47_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5994__A2 _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5861_ _3433_ _1456_ _1879_ _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7069__I _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4812_ _3461_ _0930_ _0932_ _0903_ _0933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6943__A1 _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5792_ _1029_ _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4743_ _3195_ _3139_ _0865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_109_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_30_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4674_ _0808_ _0818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6413_ _2310_ _2308_ _2420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3625_ as2650.ins_reg\[6\] _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7393_ _0204_ clknet_3_2_0_wb_clk_i as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4182__A1 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6344_ _0740_ _2352_ _2353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6857__B _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6275_ _1652_ _2273_ _2286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5226_ _1330_ _1334_ _1335_ _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6474__A3 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5157_ net5 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4108_ _0262_ _0306_ _0307_ _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5088_ _1200_ _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_38_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5434__A1 _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4237__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4039_ _3563_ _3564_ _3489_ _3573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_112_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5985__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7187__A1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_53_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6934__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_90_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6395__C1 as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3748__A1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5227__I _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4131__I _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__B _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4476__A2 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4228__A2 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3987__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_16_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6925__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3739__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4400__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4164__A1 _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4390_ as2650.holding_reg\[7\] _3248_ _0586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5900__A2 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5581__B _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4976__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3911__A1 as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7102__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6060_ _0780_ _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_input8_I io_in[7] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4467__A2 _3361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6861__B1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5011_ _0355_ _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5416__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6962_ _2382_ _2934_ _2935_ _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_53_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3978__A1 _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5913_ _1919_ _1927_ _1931_ _1932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6893_ _2219_ _2837_ _2869_ _2870_ _2227_ _2871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7332__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5844_ _1295_ _1797_ _1859_ _1863_ _1853_ _0183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A2 _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5775_ _1800_ _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6392__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4726_ _0852_ as2650.stack\[0\]\[8\] _0837_ _0853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_50_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7445_ _0256_ clknet_leaf_60_wb_clk_i as2650.psu\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6144__A2 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4657_ _0804_ _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5047__I _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3608_ as2650.cycle\[6\] _3143_ _3144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7376_ _0187_ clknet_leaf_25_wb_clk_i as2650.pc\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4588_ as2650.stack\[3\]\[0\] _0761_ _0762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6327_ _2306_ _2315_ _2336_ _2215_ _2337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6258_ _2224_ _2268_ _2269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_66_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5209_ _1237_ _1319_ _1320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6189_ _1472_ _2202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5510__I _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4630__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6907__A1 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4394__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4933__A3 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6135__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5894__A1 _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4697__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4796__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7205__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7355__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6071__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3890_ _3410_ _3417_ _3425_ _3426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3875__I as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4385__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5560_ _1597_ _1600_ _1601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_38_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_117_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4511_ _0696_ _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5491_ _1292_ _1536_ _1541_ _0152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7230_ _0041_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4442_ _0276_ _0629_ _0634_ _0010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_132_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_37_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7161_ _1349_ _1733_ _3108_ _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6200__B _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4373_ _3488_ _0569_ _0570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6112_ _2102_ _2117_ _2126_ _2127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7092_ _1137_ _3042_ _3043_ _3045_ _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_98_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6043_ _2016_ _2057_ _2058_ _2059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6854__C _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6945_ net35 _2624_ _2874_ _2921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_81_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4612__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6876_ _1553_ _0603_ _2853_ _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_74_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5827_ _1845_ _1846_ _1848_ _1849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_10_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5758_ _1695_ _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4709_ _0841_ _0838_ _0842_ _0069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6117__A2 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5689_ _0975_ _1705_ _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7428_ _0239_ clknet_leaf_2_wb_clk_i as2650.r123\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7228__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5876__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4679__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7359_ _0170_ clknet_leaf_10_wb_clk_i as2650.holding_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_78_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5891__A4 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7378__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__C _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_134_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2800 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2811 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2822 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2833 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2844 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2855 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2866 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5800__A1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2877 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2888 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2899 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_13_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_92_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7167__I _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6356__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6004__C _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6108__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5619__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6292__A1 _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4842__A2 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4991_ _1104_ _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_90_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6595__A2 _2592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6730_ _2711_ _2712_ _2670_ _2713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3942_ _3469_ _3476_ _3477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6661_ _2637_ _1807_ _1894_ _2646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6347__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3873_ _3403_ _3402_ _3408_ _3409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4358__A1 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5612_ _3207_ _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6592_ _2491_ _2590_ _2591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5543_ _1051_ _1080_ _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5570__A3 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5474_ _3207_ _1523_ _1524_ _1525_ _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_105_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5858__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7213_ _0024_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4425_ _3489_ _0600_ _0621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7144_ _1720_ _1703_ _3084_ _3095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_99_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4356_ _0541_ _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6865__B _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7075_ as2650.r123\[0\]\[6\] _3030_ _3033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4287_ _3467_ _0480_ _0484_ _0485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_140_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6283__A1 _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6026_ _2041_ _1986_ _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_80_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5060__I _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6586__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_120_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6928_ _2816_ _2903_ _2904_ _0226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_120_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6859_ _1429_ _2821_ _2838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6338__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5849__A1 _1607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5235__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5077__A2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6066__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2630 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_60 io_oeb[16] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2641 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2652 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_71 io_oeb[27] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2663 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_82 io_out[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_61_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2674 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_93 io_oeb[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__tieh
XTAP_1940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2685 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2696 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6329__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4760__A1 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6501__A2 _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5145__I _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4210_ as2650.r0\[5\] _3199_ _0409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5190_ _1161_ _3506_ _1301_ _1302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4141_ _0340_ _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5068__A2 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4072_ _3428_ _3582_ _0268_ _0272_ _0273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_96_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4974_ _3166_ _1088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5240__A2 _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_53_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6713_ _2623_ _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3925_ _3459_ _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4224__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6644_ _3187_ _2629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3856_ _3384_ _3391_ _3392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6575_ _1117_ _2505_ _2561_ _2575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3787_ _3191_ _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4200__C2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5526_ _1565_ _1569_ _1570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5457_ _3221_ _0681_ _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4408_ _0566_ _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5388_ _3181_ _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_59_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7127_ _3079_ _0250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4339_ _0438_ _0514_ _0535_ _0536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_59_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5059__A2 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7058_ _3021_ _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_41_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6009_ as2650.stack\[6\]\[2\] _1969_ _2025_ as2650.stack\[5\]\[2\] _2026_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_55_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7416__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6559__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5231__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_10_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6495__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6247__A1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6798__A2 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5470__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6970__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3710_ _3245_ _3246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_18_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3784__A2 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4690_ _0807_ _0829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3641_ _3169_ _3172_ _3174_ _3176_ _3177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_122_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6722__A2 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6360_ _2201_ _2341_ _2368_ _2369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3816__C _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4733__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5311_ as2650.r123\[3\]\[4\] _1391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6291_ _2220_ _2300_ _2301_ _2264_ _1886_ _2302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_143_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6486__A1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5242_ _1348_ _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6486__B2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5173_ _0269_ _1069_ _1285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6238__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6238__B2 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4124_ _0316_ _0317_ _0318_ _0319_ _0323_ _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_99_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7439__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6789__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput1 io_in[0] net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4219__I _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4055_ _3581_ _3588_ _3589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_83_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6862__C _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_64_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4957_ _1070_ _1071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3908_ _3442_ _3443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4888_ _3340_ _0930_ _0962_ _1004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_137_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3839_ _3374_ _3365_ _3375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6627_ _0858_ _2609_ _2613_ _0216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5516__A3 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4724__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6558_ _2013_ _0466_ _2516_ _2558_ _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5509_ _1553_ _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6489_ _3311_ _2494_ _1736_ _2495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6477__B2 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_126_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4838__B _0957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6609__I _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6229__A1 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_0_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5452__A2 _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5204__A2 _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A3 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4963__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6704__A2 _1948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5140__A1 _1202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__B1 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5860_ _1684_ _1875_ _1876_ _1878_ _1879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_62_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4811_ _3466_ _0882_ _0931_ _0932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_76_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5791_ _1814_ _1816_ _1817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_37_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4954__A1 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4742_ _0863_ _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4673_ _0710_ _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6412_ _1649_ _2230_ _2418_ _2419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3624_ _3159_ _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4706__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7392_ _0203_ clknet_leaf_9_wb_clk_i as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6343_ _0734_ _2317_ _2352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4182__A2 _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__C _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6274_ _1903_ _2284_ _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_131_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7261__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5225_ _1130_ _1329_ _1335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5131__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5682__A2 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5156_ _0609_ _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4107_ as2650.holding_reg\[3\] _3258_ _0307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5087_ _0863_ _3236_ _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_72_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5434__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6631__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4038_ _3444_ _3571_ _3488_ _3572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_84_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3788__I _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7187__A2 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__B1 _2027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5989_ _2003_ _2004_ _2005_ _2006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XPHY_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__C2 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3748__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6147__B1 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5508__I _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6767__C _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3920__A2 _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6870__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3684__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5399__B _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3987__A2 _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5189__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_43_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6023__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6689__A1 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7284__CLK clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_27_wb_clk_i_I clknet_opt_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_3_4_0_wb_clk_i clknet_0_wb_clk_i clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_67_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A1 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5010_ _3179_ _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6861__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6861__B2 _2839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5416__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6613__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6961_ _2934_ _2935_ _2382_ _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_53_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5912_ _1473_ _1928_ _1930_ _1931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3978__A2 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6892_ _1428_ _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_74_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_34_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5843_ _1179_ _1861_ _1862_ _1863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_61_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5719__A3 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4927__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5774_ _1799_ _1800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4725_ _0730_ _0852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7444_ _0255_ clknet_leaf_52_wb_clk_i net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4656_ _0779_ as2650.stack_ptr\[0\] _0804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3607_ _3141_ _3142_ _3143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5352__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4587_ _0758_ _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7375_ _0186_ clknet_leaf_47_wb_clk_i as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6326_ _2314_ _2327_ _2335_ _2336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5104__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6257_ as2650.pc\[7\] _1211_ _2180_ _2267_ _2268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_118_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6852__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5208_ _1318_ _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6188_ _1742_ _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_112_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6095__S _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5139_ _1205_ _1245_ _1251_ _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_123_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6604__A1 as2650.stack\[7\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_8_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_8_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4407__I _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4091__A1 _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6907__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4142__I _0341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_126_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5894__A2 _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A1 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7121__C _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4317__I _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4082__A1 _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4909__A1 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5582__A1 _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4510_ _0695_ _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5490_ _1540_ _1538_ _1541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4441_ as2650.r123\[1\]\[2\] _0631_ _0634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5334__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4987__I _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5885__A2 _1902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7160_ _3107_ _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4372_ _0568_ _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6111_ _1818_ _2094_ _2125_ _2088_ _2126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7091_ _1566_ _1066_ _1179_ _1173_ _3044_ _3045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6834__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6042_ _3538_ _2014_ _2058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5611__I _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6944_ _2304_ _2788_ _2913_ _2916_ _2919_ _2920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_82_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_23_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_41_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5767__B _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6875_ _2851_ _2830_ _2852_ _2853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6442__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5826_ _3184_ _3314_ _1847_ _1619_ _1848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_23_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4376__A2 _0435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A1 _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5757_ _1436_ _1775_ _1777_ _1778_ _1783_ _1784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_4708_ as2650.stack\[0\]\[1\] _0839_ _0842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6117__A3 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5688_ _1720_ _1641_ _1721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7427_ _0238_ clknet_leaf_14_wb_clk_i net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5325__A1 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4128__A2 as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6522__B1 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4639_ _0718_ _0791_ _0794_ _0047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7358_ _0169_ clknet_3_0_0_wb_clk_i as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7078__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6309_ _2007_ _2312_ _2319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7289_ _0100_ clknet_leaf_50_wb_clk_i as2650.stack\[6\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_133_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4300__A2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2801 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2812 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6053__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2823 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2834 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2845 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2856 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2867 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2878 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2889 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7002__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5564__A1 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7322__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5619__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6292__A2 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4990_ _0357_ _1104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3941_ _3472_ _3475_ _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6660_ _1134_ _1511_ _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3872_ _3407_ _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5611_ _1134_ _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4358__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6591_ _1351_ _1264_ _1265_ _2589_ _1516_ _2590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_129_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5542_ _1145_ _1167_ _1163_ _1518_ _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_117_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_9_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__B1 _2507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5473_ _0680_ _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5858__A2 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4424_ _3444_ _0603_ _0616_ _0619_ _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7212_ _0023_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3869__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7143_ _3432_ _3093_ _3094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4355_ _0551_ _0543_ _0552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6807__A1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7074_ _0510_ _3029_ _3032_ _0244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4286_ _0483_ _3469_ _3371_ _0484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6025_ as2650.pc\[3\] _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6035__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6927_ net50 _2786_ _2874_ _2904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5794__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6858_ _2648_ _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5809_ _1695_ _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5546__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6789_ _2763_ _0330_ _2770_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_104_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6274__A2 _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5251__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6026__A2 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2620 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2631 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A1 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2642 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_61 io_oeb[17] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2653 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_72 io_oeb[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_83 io_out[28] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2664 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4588__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2675 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2686 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2697 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4760__A2 _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4140_ _0335_ _0339_ _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_123_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5068__A3 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4071_ _3419_ _0271_ _3397_ _0272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4276__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4973_ _1081_ _1084_ _1086_ _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_6712_ _2625_ _2693_ _2695_ _0219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4505__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3924_ _3458_ _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_75_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6643_ _2627_ _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3855_ _3390_ _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3786_ _3137_ _3321_ _3322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4200__A1 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6574_ _2541_ _0537_ _2542_ _2573_ _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4200__B2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5525_ _1567_ _1166_ _1164_ _1568_ _1569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5456_ _1133_ _1506_ _1430_ _1507_ _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_86_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4407_ _0602_ _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5700__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5387_ _0356_ _1133_ _0673_ _1449_ _1450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_132_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7126_ _1736_ _3077_ _3078_ _3079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_82_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4338_ _0530_ _0534_ _0535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7057_ _3288_ _1042_ _3021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4269_ _0466_ _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_75_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4267__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6008_ _1970_ _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A1 _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4415__I _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5519__A1 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6495__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_133_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4258__A1 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6540__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3640_ _3175_ _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6183__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5156__I _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5310_ _1390_ _0122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6290_ _2176_ _2275_ _2184_ _2301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6486__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5241_ _1214_ _1348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_102_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5172_ _1043_ _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6238__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4123_ _0320_ _0321_ _0322_ _0323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_122_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xinput2 io_in[1] net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4054_ _3500_ _3583_ _3508_ _3587_ _3588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_84_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6410__A2 _2373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7190__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4956_ _3327_ _1069_ _1062_ _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3907_ _3188_ _3277_ _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_138_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4887_ _0559_ _0978_ _0889_ _1002_ _1003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_137_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6626_ as2650.stack\[7\]\[11\] _2610_ _2613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3838_ _3373_ _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5516__A4 _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_14_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6557_ _1764_ _0475_ _2557_ _2499_ _2558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3769_ _3143_ _3304_ _3183_ _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_118_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5508_ _1014_ _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6488_ _2490_ _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_10_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6477__A2 _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5439_ _1127_ _1490_ _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_133_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7109_ _3500_ _3523_ _0273_ _3061_ _3062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_59_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5988__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output22_I net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4145__I _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6401__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5755__A4 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5685__B _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4963__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5912__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_17_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7114__B1 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6468__A2 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4479__A1 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5140__A2 _1252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5979__B2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4651__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4810_ _3476_ _0886_ _0887_ _0931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5790_ _1815_ _1635_ _1816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA_clkbuf_leaf_56_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4741_ _0862_ _0863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4954__A2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4672_ _0815_ _0809_ _0816_ _0058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6411_ _0747_ _2417_ _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3623_ as2650.ins_reg\[5\] _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4706__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7391_ _0202_ clknet_leaf_10_wb_clk_i as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_127_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6342_ _1542_ _2350_ _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4939__B _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7406__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6273_ _1891_ _1453_ _2284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5224_ _1333_ _1319_ _1334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5131__A2 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5155_ as2650.r0\[7\] _1266_ _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4890__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4106_ _0282_ _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5086_ _3414_ _3508_ _0295_ _1192_ _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_84_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4037_ _3566_ _3570_ _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_112_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A1 as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5988_ _1240_ _2004_ _2005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_36_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4939_ _0678_ _1045_ _1052_ _1053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_21_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6147__B2 as2650.stack\[5\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6609_ _2594_ _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_opt_1_0_wb_clk_i clknet_3_3_0_wb_clk_i clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_10_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5524__I _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6870__A2 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4881__A1 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6622__A2 _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4633__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5189__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6304__B _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6138__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7429__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6689__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6958__C _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6974__B _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6861__A2 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6265__I as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6613__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6960_ _2308_ _2895_ _2935_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_93_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5672__I0 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5911_ as2650.stack\[7\]\[0\] _1929_ _1925_ as2650.stack\[6\]\[0\] _1930_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6891_ _2235_ _2868_ _2869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_46_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5842_ _1071_ _1267_ _3237_ _1862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5719__A4 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5773_ _1143_ _1589_ _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5609__I _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6129__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4724_ _0850_ _0845_ _0851_ _0075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7443_ _0254_ clknet_3_4_0_wb_clk_i as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4655_ _0749_ _0798_ _0803_ _0054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3606_ as2650.cycle\[5\] as2650.cycle\[4\] _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7374_ _0185_ clknet_3_5_0_wb_clk_i as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5352__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4586_ _0759_ _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6325_ _2201_ _2306_ _2334_ _2335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5344__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6256_ _2177_ _2223_ _2267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5104__A2 _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5207_ _1317_ _3304_ _1318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6852__A2 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6187_ _1812_ _2199_ _2200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_57_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4863__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5138_ _1138_ _1208_ _1248_ _1250_ _1251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_85_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6604__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5069_ _1137_ _1148_ _1159_ _1181_ _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4615__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5591__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7096__A2 _3049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6843__A2 _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3901__I0 _3394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7251__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4909__A2 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5429__I _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4440_ _3526_ _0629_ _0633_ _0009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6531__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4371_ _0316_ _0566_ _0540_ _0319_ _0567_ _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_98_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6110_ _1030_ _2120_ _2124_ _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7087__A2 _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7090_ _1579_ _1250_ _3044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6041_ _3538_ _2014_ _2057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4845__A1 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_47_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_47_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_67_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6943_ _2313_ _2918_ _2919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6874_ _1272_ _0546_ _2852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5825_ _1831_ _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5022__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5756_ _1779_ _1782_ _1783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6770__A1 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5783__B _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4707_ _0696_ _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5687_ _1719_ _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7426_ _0237_ clknet_leaf_15_wb_clk_i net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6522__A1 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5325__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4638_ as2650.stack\[2\]\[5\] _0792_ _0794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6522__B2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7357_ _0168_ clknet_leaf_65_wb_clk_i as2650.holding_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4569_ _0744_ _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6308_ _2304_ _2317_ _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7288_ _0099_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5089__B2 _1199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6239_ as2650.stack\[6\]\[7\] _1925_ _2030_ _2251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4836__A1 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6589__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2802 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2813 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7274__CLK clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2824 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2835 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2846 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2857 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2868 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2879 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7002__A2 _2973_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5249__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5693__B _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5619__A3 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6808__I _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5868__B _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5252__A1 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3940_ _3369_ _3473_ _3474_ _3475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_90_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3871_ _3404_ _3406_ _3407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5610_ _1146_ _1649_ _1609_ _1650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5555__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6590_ _1295_ _1092_ _2588_ _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4358__A3 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6699__B _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5541_ _1516_ _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_125_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5960__C1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5472_ _0679_ _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6504__B2 _2508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7211_ _0022_ clknet_leaf_36_wb_clk_i as2650.stack\[4\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4423_ _0618_ _0359_ _0361_ _0619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5858__A3 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7142_ _3088_ _3092_ _3093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4354_ _3282_ _0396_ _0372_ _0449_ _0551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_141_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6718__I _1676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7073_ as2650.r123\[0\]\[5\] _3030_ _3032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_101_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4285_ _0482_ _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4818__A1 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6024_ _0702_ _1984_ _2040_ _0186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7297__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5491__A1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5778__B _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4046__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5243__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6453__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6926_ _0730_ _2788_ _2897_ _2692_ _2902_ _2903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_54_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6857_ _1832_ _2819_ _2835_ _2455_ _2836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
Xfanout46 net48 net46 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_23_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5808_ _1553_ _1637_ _1833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5546__A2 _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6788_ _1719_ _2629_ _2667_ _2768_ _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_52_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5739_ _1307_ _1636_ _1766_ _1767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_109_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7409_ _0220_ clknet_opt_3_1_wb_clk_i net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2610 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2621 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2632 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4037__A2 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2643 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__B1 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_62 io_oeb[18] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2654 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_73 io_oeb[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2665 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_84 io_out[29] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2676 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2687 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2698 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5537__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5707__I _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4760__A3 _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5170__B1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4070_ _0269_ _3579_ _0270_ _0271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_84_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4276__A2 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_97_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3897__I _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A1 _1130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4972_ _1085_ _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6973__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6711_ net52 _2654_ _2694_ _2695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3923_ _3455_ _3457_ _3458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6642_ _1503_ _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3854_ _3297_ _3389_ _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6725__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6573_ _2447_ _2571_ _2572_ _2573_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_118_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3785_ as2650.r123\[2\]\[7\] as2650.r123_2\[2\]\[7\] _3193_ _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_118_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4521__I _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5524_ _1444_ _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5455_ _3271_ _1449_ _1507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_117_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7150__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_62_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4406_ _3339_ _3389_ _0599_ _3567_ _0601_ _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5161__B1 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5386_ _0660_ _1448_ _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5700__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7125_ _3050_ _3075_ _3411_ _3078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4337_ _3423_ _0532_ _0533_ _0279_ _0534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_119_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7056_ _3002_ _3019_ _3020_ _0238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4268_ _0438_ _0462_ _0464_ _0465_ _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_87_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_101_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4267__A2 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6007_ _1472_ _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4199_ _0340_ _0321_ _0398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_70_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6964__A1 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A2 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6909_ _0610_ _0622_ _2886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5519__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3950__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7141__A1 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5455__A1 _3271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4258__A2 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5207__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6955__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_46_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4430__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6707__A1 _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6707__B2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5437__I _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5881__B _1899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3941__A1 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5240_ _1330_ _1346_ _1347_ _0095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4497__A2 _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5171_ _3253_ _0424_ _1278_ _1282_ _1283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_64_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4122_ _3459_ _3553_ _0306_ _0322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_111_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4053_ _3585_ _3402_ _3586_ _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_83_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput3 io_in[2] net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_83_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4516__I _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7335__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6946__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4955_ _1068_ _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3906_ _3290_ _3437_ _3441_ _0000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4886_ _0556_ _0977_ _1002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_32_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7048__B _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6625_ _0740_ _2609_ _2612_ _0215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3837_ _3372_ _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4251__I _0448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6556_ _1519_ _0505_ _2557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_3768_ _3182_ _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5507_ _1236_ _1547_ _1552_ _0157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_3_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7123__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6487_ _2454_ _2456_ _2467_ _1583_ _2492_ _2493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3699_ _3140_ _3234_ _3235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5438_ _1489_ _1419_ _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5685__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6178__I _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5369_ _3169_ _3151_ _0672_ _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_120_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7108_ _0901_ _3460_ _3060_ _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7039_ net40 _3000_ _3008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6937__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output15_I net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4412__A2 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4963__A3 _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3923__A1 _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7114__B2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7208__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4479__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A1 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7358__CLK clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5979__A2 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_2_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6928__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4403__A2 _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4740_ _3254_ _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4954__A3 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4671_ as2650.stack\[1\]\[3\] _0810_ _0816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5167__I as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6156__A2 _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6410_ _2413_ _2373_ _2352_ _2417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4167__A1 _3290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3622_ as2650.ins_reg\[4\] _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7390_ _0201_ clknet_leaf_9_wb_clk_i as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6341_ _2276_ _2349_ _1744_ _2278_ _2350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_116_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__A1 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6272_ _0729_ _2282_ _2283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_100_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5223_ _1238_ _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5131__A3 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_130_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5154_ _1249_ _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4105_ _3404_ _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_99_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5085_ _1183_ _1197_ _1198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6092__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4036_ _3567_ _3568_ _3569_ _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_112_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6919__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5987_ _1452_ _2004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6395__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_52_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4938_ _1049_ _1051_ _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1002 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4869_ _0974_ _0944_ _0986_ _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6147__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4158__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6608_ _2595_ _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6539_ _2446_ _2541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4849__C _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4330__A1 as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3684__A3 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4881__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_60_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5830__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4633__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4156__I _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_71_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3995__I _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6304__C _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6138__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4149__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5897__A1 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5649__A1 _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6310__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5113__A3 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6974__C _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_87_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_66_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5821__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5672__I1 _1707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5910_ _0649_ _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6890_ _1745_ _2860_ _2868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_4_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5841_ _1295_ _1351_ _1860_ _1861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_22_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4388__A1 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5772_ _1575_ _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_21_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4723_ as2650.stack\[0\]\[7\] _0846_ _0851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7442_ _0253_ clknet_leaf_54_wb_clk_i as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4654_ as2650.stack\[2\]\[12\] _0799_ _0803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5888__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3605_ as2650.cycle\[7\] _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7373_ _0184_ clknet_leaf_25_wb_clk_i as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4585_ _0758_ _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6324_ _2202_ _2330_ _2333_ _2211_ _2334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4560__A1 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6255_ _2265_ _2266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_89_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5104__A3 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5206_ _3147_ _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6186_ _2190_ _2192_ _2198_ _2065_ _2199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_112_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__A2 _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5137_ _1143_ _1249_ _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5360__I _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6065__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5068_ _1172_ _1176_ _1177_ _1180_ _1181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_72_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4019_ _3552_ _3553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_25_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_52_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_80_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4379__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4704__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5591__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__C _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5535__I _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3901__I1 _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6056__B2 _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__B1 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4790__A1 _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4370_ _3574_ _0542_ _0567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_125_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7087__A3 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6040_ _1453_ _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input6_I io_in[5] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5180__I _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6047__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6942_ _2304_ _2837_ _2917_ _2870_ _1939_ _2918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_82_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_16_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_16_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_6873_ _1213_ _0545_ _2851_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_23_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5824_ _1823_ _1844_ _1675_ _1846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5022__A2 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5755_ _1781_ _1490_ _1649_ _1778_ _1782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_124_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6770__A2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5573__A3 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5783__C _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4781__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4706_ _0835_ _0838_ _0840_ _0068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5686_ _1289_ _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7425_ _0236_ clknet_leaf_15_wb_clk_i net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4637_ _0711_ _0791_ _0793_ _0046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5355__I _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6522__A2 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4568_ _0743_ _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7356_ _0167_ clknet_leaf_65_wb_clk_i as2650.holding_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6307_ _0728_ _2219_ _2231_ _2317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_103_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7287_ _0098_ clknet_leaf_49_wb_clk_i as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4499_ _0683_ _3274_ _0685_ _0686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5291__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5089__A2 _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6286__A1 _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6238_ as2650.stack\[5\]\[7\] _2025_ _2027_ as2650.stack\[4\]\[7\] as2650.stack\[7\]\[7\]
+ _0650_ _2250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_103_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6169_ _2178_ _2181_ _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5090__I _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_40_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2803 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2814 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2825 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2836 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2847 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2858 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2869 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4434__I _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6277__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5619__A4 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_27_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4609__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6029__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5252__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3870_ _3405_ _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5540_ net20 _1582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4763__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__B1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5960__C2 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5471_ _3362_ _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_69_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6504__A2 _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7210_ _0021_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4422_ _0617_ _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_67_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7141_ _1076_ _1118_ _1086_ _3091_ _3092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
X_4353_ _3340_ _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5903__I _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6268__A1 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7072_ _0434_ _3029_ _3031_ _0243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4284_ _0481_ _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_141_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6023_ _1985_ _2038_ _2039_ _2040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5243__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6925_ _2220_ _2901_ _2902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6856_ _2638_ _2821_ _2834_ _1828_ _2835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_39_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xfanout47 net48 net47 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_22_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5807_ _1831_ _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_56_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3999_ as2650.r123\[0\]\[3\] as2650.r123\[2\]\[3\] as2650.r123_2\[0\]\[3\] as2650.r123_2\[2\]\[3\]
+ _3196_ _3349_ _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__5286__S _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6787_ _2629_ _2767_ _2768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4754__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5738_ _1527_ _1676_ _1766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_136_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6402__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5669_ _1097_ _1705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7408_ _0219_ clknet_leaf_27_wb_clk_i net26 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7339_ _0150_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7241__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A2 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output45_I net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6644__I _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2600 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2611 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2622 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2633 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A1 as2650.stack\[3\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2644 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_63 io_oeb[19] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_3389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_36_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_74 io_oeb[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_2_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2655 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2666 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_85 io_out[30] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XANTENNA__6982__A2 _2936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2677 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2688 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2699 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4993__A1 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__B1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5537__A3 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6498__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5170__A1 _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5170__B2 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6670__A1 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5225__A2 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4971_ _0336_ _1068_ _1062_ _1085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_63_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6973__A2 _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6710_ _1459_ _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3922_ _3198_ _3456_ _3457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4984__A1 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6641_ _1498_ _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3853_ _3386_ _3388_ _3389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_4
XFILLER_20_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4736__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3784_ as2650.r0\[7\] _3199_ _3320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6572_ _2452_ _0569_ _2572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_125_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5523_ _1566_ _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_121_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6489__A1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5454_ _0670_ _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7150__A2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7264__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4405_ _3565_ _0600_ _0601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5161__A1 _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5385_ _3266_ _0656_ _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5161__B2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4336_ _0531_ _0497_ _3517_ _0533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7124_ _3056_ _3057_ _3074_ _3076_ _3077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7055_ net44 _2992_ _3020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4267_ _0438_ _0439_ _0465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6661__A1 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6006_ _1999_ _2022_ _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_31_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4198_ _0396_ _0341_ _0397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_91_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5767__A3 _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6908_ _2845_ _2824_ _2884_ _2846_ _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_4
XFILLER_70_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6839_ _2180_ _2817_ _2818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_50_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5455__A2 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5207__A2 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3769__A2 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4966__A1 _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6323__B _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7287__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A1 _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5881__C _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4497__A3 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6891__A1 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5170_ _1279_ _3464_ _1280_ _1117_ _1281_ _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_96_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4121_ _0263_ _3552_ _0283_ _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_110_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4052_ _3421_ _3427_ _3586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_111_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xinput4 io_in[3] net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XANTENNA__5402__B _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3701__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4406__B1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4954_ _3179_ _3173_ _3356_ _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3905_ as2650.r123\[2\]\[0\] _3440_ _3441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_71_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4885_ _0864_ _3272_ _0865_ _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__4709__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6624_ as2650.stack\[7\]\[10\] _2610_ _2612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3836_ net1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5382__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6555_ _2546_ _2554_ _2556_ _0201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3767_ _3255_ _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5506_ _3229_ _1549_ _1552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_134_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6486_ _3370_ _1524_ _1850_ _3548_ _2491_ _2492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3698_ _3190_ _3201_ _3223_ _3233_ _3234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_118_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5134__A1 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5437_ _0660_ _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5363__I _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5685__A2 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5368_ _1430_ _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7107_ _0261_ _0901_ _3060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4319_ _0447_ _0459_ _0373_ _0385_ _0440_ _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_101_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5299_ _1384_ _1375_ _1385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A1 _1526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7038_ _0354_ _2996_ _3006_ _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_75_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4707__I _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6937__A2 _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4948__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5966__C _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_71_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4963__A4 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6797__C _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6322__B1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5273__I _1353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5676__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3687__A1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6625__A1 _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7050__A1 _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4553__S _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4352__I _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4670_ _0705_ _0815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__B _1906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3621_ _3156_ _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4167__A2 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6340_ _2321_ _2349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_127_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7105__A2 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6271_ _2219_ _2231_ _2282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6864__A1 _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5222_ _1320_ _1330_ _1332_ _0092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_116_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5153_ _1223_ _0613_ _1221_ _1263_ _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__7302__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4104_ _3261_ _3536_ _0302_ _0303_ _0304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_96_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5084_ _1188_ _1195_ _1196_ _1197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4527__I _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6092__A2 _2100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4035_ _3388_ _3460_ _3565_ _3569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_38_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_129_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5986_ as2650.addr_buff\[2\] _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_53_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_75_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7059__B _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4937_ _1050_ _1028_ _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4262__I _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4868_ _0400_ _0908_ _0985_ _0910_ _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6607_ _0705_ _2596_ _2601_ _0208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3819_ _3354_ _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4799_ _3432_ _3140_ _3265_ _0920_ _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_134_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3905__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6538_ _2539_ _2540_ _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_106_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6469_ _2471_ _2473_ _2474_ _2475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3669__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6607__A1 _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4094__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5830__A2 _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5346__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5897__A2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7099__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5217__B _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7099__B2 _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7325__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6846__A1 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5649__A2 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_78_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6074__A2 _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7023__A1 _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5840_ _1130_ _1351_ _1860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_35_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5771_ _1774_ _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5178__I net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4722_ _0725_ _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7441_ _0252_ clknet_leaf_60_wb_clk_i as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_2
XANTENNA__5337__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6534__B1 _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4653_ _0745_ _0798_ _0802_ _0053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5906__I _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3604_ _3139_ _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5888__A2 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7372_ _0183_ clknet_leaf_52_wb_clk_i as2650.psu\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__A1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4584_ _0755_ _0757_ _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6323_ _2331_ _2332_ _2209_ _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6254_ as2650.pc\[8\] _0558_ _2265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5205_ _1255_ _1182_ _1316_ _1116_ _0091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4312__A2 _0467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6185_ _2066_ _2193_ _2196_ _2197_ _2198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_69_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5136_ _3152_ _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_44_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5067_ _1173_ _1179_ _1180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_84_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5797__B _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4018_ _3135_ _3550_ _3551_ _3295_ _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_72_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5289__S _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7014__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6405__C _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5576__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4379__A2 _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5969_ as2650.pc\[2\] _1937_ as2650.pc\[0\] _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__5088__I _1200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5591__A4 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5328__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7348__CLK clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4000__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A1 _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4303__A2 _0500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7005__A1 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5567__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5567__B2 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1075 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4542__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5461__I _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6047__A2 _2062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4058__A1 _3591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6941_ _2151_ _2906_ _2322_ _2917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3805__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4805__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6872_ _2662_ _2848_ _2849_ _2628_ _2850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5823_ _1675_ _1823_ _1844_ _1845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5558__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5754_ _1780_ _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_56_wb_clk_i clknet_3_4_0_wb_clk_i clknet_leaf_56_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5573__A4 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4705_ as2650.stack\[0\]\[0\] _0839_ _0840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6507__B1 _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5685_ _0281_ _1709_ _1718_ _0169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4540__I _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7424_ _0235_ clknet_leaf_15_wb_clk_i net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4636_ as2650.stack\[2\]\[4\] _0792_ _0793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7355_ _0166_ clknet_leaf_65_wb_clk_i as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5730__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4567_ as2650.pc\[11\] _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_143_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6306_ _1540_ _2280_ _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7286_ _0097_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4498_ _0684_ _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_104_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6237_ _2064_ _2241_ _2248_ _2249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_77_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5371__I _0668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4297__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6168_ _2136_ _2134_ _2180_ _2181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5119_ _0884_ _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6099_ _1289_ _1806_ _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_58_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2804 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5797__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2815 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2826 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2837 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2848 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4715__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2859 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_3_0_wb_clk_i clknet_0_wb_clk_i clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XANTENNA__6135__C _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5549__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4524__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6277__A2 _2285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_65_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5788__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4625__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4763__A2 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5960__A1 as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4360__I net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5470_ _1075_ _1511_ _1515_ _1521_ _1522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__6996__B as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4421_ as2650.r0\[7\] _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5712__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7140_ _1056_ _1108_ _3090_ _3091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4352_ _0463_ _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4283_ net6 _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7071_ as2650.r123\[0\]\[4\] _3030_ _3031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_99_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6022_ _1469_ _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5779__A1 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5140__B _1182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6924_ _0729_ _2721_ _2900_ _2720_ _2901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_70_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6855_ _2827_ _2833_ _2747_ _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xfanout48 net49 net48 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5806_ _1766_ _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6786_ _0424_ _0400_ _2766_ _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_50_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_3998_ _3132_ _3530_ _3531_ _3332_ _3532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5737_ _1761_ _1762_ _1764_ _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5366__I _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5668_ _1333_ _1703_ _1704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7407_ _0218_ clknet_leaf_27_wb_clk_i net25 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4619_ _0779_ _0751_ _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5599_ _1639_ _1156_ net49 _1640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_2_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7338_ _0149_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_137_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7269_ _0080_ clknet_leaf_32_wb_clk_i as2650.stack\[0\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2601 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__B1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2612 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output38_I net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4445__I _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2623 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2634 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6431__A2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xwrapped_as2650_53 io_oeb[9] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2645 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_64 io_oeb[20] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2656 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_75 io_oeb[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2667 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_86 io_out[31] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2678 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2689 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A2 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_9_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6195__B2 as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5942__A1 _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4180__I _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_1_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6498__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5170__A2 _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6670__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4783__C _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6422__A2 _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4970_ _1082_ _1083_ _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3921_ as2650.r123\[0\]\[2\] as2650.r123\[2\]\[2\] as2650.r123_2\[0\]\[2\] as2650.r123_2\[2\]\[2\]
+ _3131_ _3349_ _3456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__4984__A2 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6640_ _2624_ _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6186__A1 _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3852_ as2650.addr_buff\[5\] _3387_ _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6186__B2 _2065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6503__C _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6571_ _2450_ _0546_ _2571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5933__A1 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3783_ as2650.psl\[3\] _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5522_ _0896_ _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_121_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6489__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5453_ _1491_ _1504_ _1200_ _1505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7150__A3 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4404_ _3337_ _0538_ _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5161__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5384_ _1438_ _1446_ _1447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_99_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7123_ _3050_ _3075_ _3076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4335_ _0531_ _0497_ _0532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_59_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7054_ _2991_ _2577_ _3018_ _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6110__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4266_ _0458_ _0312_ _0463_ _0464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_86_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6005_ _2000_ _2012_ _2021_ _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_86_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6661__A2 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_41_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4197_ _0395_ _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_83_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6413__A2 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4265__I _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6907_ _0609_ _0622_ _2884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4975__A2 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6838_ _2133_ _2789_ _2817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6177__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5924__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6769_ _1242_ _2191_ _2751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_10_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7141__A3 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6655__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A2 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_34_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4966__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4718__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5391__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4120_ as2650.idx_ctrl\[1\] _3186_ _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4051_ _3584_ as2650.carry _3585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_68_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4654__A1 as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput5 io_in[4] net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_83_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_25_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4406__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4018__C _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4953_ _0893_ _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_33_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3904_ _3439_ _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_36_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6159__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4884_ _1000_ _0086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6623_ _0734_ _2609_ _2611_ _0214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_20_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3835_ _3344_ _3371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4709__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6554_ _0975_ _2555_ _2217_ _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3766_ _3301_ _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5382__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3873__B _3408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5505_ _1235_ _1547_ _1551_ _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6485_ _2490_ _2491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3697_ _3205_ _3227_ _3232_ _3233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_133_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5436_ _1291_ _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_133_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6331__A1 as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5134__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_138_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_3_1_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5367_ _0681_ _1430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_47_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4893__A1 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7106_ _3500_ _3522_ _3421_ _3430_ _3059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4318_ _0458_ _0460_ _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5298_ _1011_ _1384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_87_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7037_ _2997_ _0976_ _3006_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4249_ as2650.holding_reg\[5\] _0447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_87_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_27_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6398__B2 _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6570__A1 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6322__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6873__A2 _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6625__A2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3802__I _3337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4636__A1 as2650.stack\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7254__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4939__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5665__S _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6988__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3620_ _3155_ _3156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6561__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5364__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6270_ _2276_ _2279_ _2280_ _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6313__A1 _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5221_ _1061_ _1331_ _1332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6864__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4875__A1 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5152_ _1263_ _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4103_ _3406_ _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_69_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6616__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4808__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5083_ _0579_ _0582_ _1188_ _1195_ _1196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_42_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4034_ _3545_ _3553_ _3568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_65_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3850__A2 as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5985_ _0700_ _2001_ _2002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5052__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4936_ _3357_ _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4867_ _0947_ _0983_ _0984_ _0985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6606_ as2650.stack\[7\]\[3\] _2597_ _2601_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_123_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3818_ _3353_ _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6552__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4798_ _0919_ _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6537_ _0354_ _2494_ _1461_ _2540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3749_ _3284_ _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_115_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6468_ _3265_ _0920_ _1152_ _1158_ _2474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5419_ _1478_ _0143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6399_ _2398_ _2399_ _2406_ _2407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_121_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4866__A1 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3669__A2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6607__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3622__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7277__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4094__A2 _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_55_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_43_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5043__A1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5346__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7099__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6846__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4306__B1 _0469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_opt_1_0_wb_clk_i_I clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5459__I _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5770_ _1773_ _1796_ _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5585__A2 _1625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4721_ _0823_ _0845_ _0849_ _0074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7440_ _0251_ clknet_leaf_6_wb_clk_i as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6534__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4652_ as2650.stack\[2\]\[11\] _0799_ _0802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3603_ as2650.halted net10 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7371_ _0182_ clknet_3_3_0_wb_clk_i as2650.cycle\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_50_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4583_ _0652_ _0756_ _0757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3899__A2 _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6322_ as2650.stack\[3\]\[9\] _0649_ _0781_ as2650.stack\[1\]\[9\] _2332_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_143_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6253_ _0729_ _2263_ _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_48_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4848__A1 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5204_ _1182_ _1315_ _1316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6184_ _1348_ _1513_ _1815_ _3229_ _1210_ _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__6239__B _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5135_ _0598_ _1247_ _1248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_111_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5066_ _1060_ _1178_ _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_38_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_16_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4076__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4017_ _3346_ _3347_ _3551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5797__C _1822_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5025__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6773__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5968_ _1882_ _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6773__B2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4919_ _1032_ _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5899_ _1151_ _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6525__A1 _2527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5328__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4000__A2 _3533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__A2 _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4892__B _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A1 as2650.stack\[6\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5016__A1 _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5567__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6764__A1 _1544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5319__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7442__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4058__A2 _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5255__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_54_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6940_ _2861_ _2915_ _2866_ _2916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_47_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3805__A2 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6871_ _1231_ _2662_ _2849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5007__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5822_ as2650.cycle\[5\] _1839_ _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6755__A1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5558__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5753_ _1084_ _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4230__A2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5917__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4704_ _0836_ _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6507__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5684_ _1700_ _1716_ _1717_ _1718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7423_ _0234_ clknet_leaf_15_wb_clk_i net40 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_136_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4635_ _0783_ _0792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7354_ _0165_ clknet_leaf_12_wb_clk_i as2650.idx_ctrl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
Xclkbuf_leaf_25_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4566_ _0741_ _0736_ _0742_ _0026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6305_ _2176_ _2314_ _2184_ _2315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3741__A1 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7285_ _0096_ clknet_leaf_8_wb_clk_i as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4497_ _3267_ _3216_ _3213_ _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_131_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6236_ _1307_ _2013_ _2245_ _2247_ _2053_ _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XANTENNA__5494__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6167_ _0716_ _0482_ _2179_ _2180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5118_ _0611_ _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_3506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6098_ _1289_ _2110_ _2112_ _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XTAP_3517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4049__A2 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5246__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5049_ _1161_ _1154_ _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XTAP_2805 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3900__I _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2816 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6994__A1 net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5797__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2827 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2838 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2849 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5099__I _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6746__A1 _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5549__A2 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A2 _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__B1 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_4_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3810__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6985__A1 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5788__A2 _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3799__A1 _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5938__S _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A1 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5960__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7162__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4420_ _3450_ _0604_ _0615_ _3313_ _0616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5712__A2 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4351_ _0547_ _0359_ _0548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5472__I _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7070_ _3023_ _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4282_ _0460_ _0479_ _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_113_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6021_ _1988_ _1998_ _2036_ _2037_ _2038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA_clkbuf_3_6_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4816__I _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7338__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A2 _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3720__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6236__C _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6923_ _2000_ _2286_ _2898_ _2899_ _2900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_39_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6854_ _2671_ _2831_ _2832_ _2448_ _2833_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_62_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xfanout49 net18 net49 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
X_5805_ _1762_ _1825_ _1829_ _1830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_50_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_56_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6785_ _2764_ _2765_ _2766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3997_ as2650.r0\[3\] _3331_ _3531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5400__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4551__I _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5736_ _1763_ _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_52_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4754__A3 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7153__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5667_ _1149_ _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5164__B1 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4618_ as2650.stack_ptr\[1\] _0779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7406_ _0217_ clknet_leaf_33_wb_clk_i as2650.stack\[7\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5598_ _1431_ _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7337_ _0148_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4549_ as2650.pc\[8\] _0728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7268_ _0079_ clknet_leaf_37_wb_clk_i as2650.stack\[0\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6664__B1 _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6219_ _0721_ _2142_ _2231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_77_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7199_ _0010_ clknet_leaf_1_wb_clk_i as2650.r123\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_63_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5482__A4 _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A1 _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6427__B _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__A1 _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2602 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6967__B2 _2941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2613 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2624 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2635 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_54 io_oeb[10] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_65 io_oeb[21] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_2646 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4442__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2657 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_76 io_oeb[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2668 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_87 io_out[32] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_60_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2679 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6719__A1 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4993__A3 _1106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6195__A2 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7144__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6958__A1 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6422__A3 _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5630__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4433__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3920_ _3132_ _3453_ _3454_ _3332_ _3455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_44_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7168__B _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3851_ as2650.addr_buff\[6\] _3387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6186__A2 _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6570_ _2494_ _2568_ _2570_ _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3782_ _3317_ _3318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4304__C _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5933__A2 _1950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5521_ _1448_ _1129_ _1565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_74_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7135__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5452_ _1494_ _1499_ _1503_ _1504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_51_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4403_ _3338_ _0598_ _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_126_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5383_ _1439_ _1266_ _1442_ _1445_ _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_126_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7122_ _1237_ _1692_ _1150_ _3075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4334_ as2650.holding_reg\[6\] _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5449__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7053_ _0618_ _2997_ _3018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4265_ _0460_ _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6004_ _2013_ _2017_ _2018_ _2020_ _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4121__A1 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4196_ _3296_ _3470_ _0263_ _0283_ _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__6247__B _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4672__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4546__I _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6949__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4424__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6906_ _1537_ _2882_ _2883_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_93_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6837_ _2726_ _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_11_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6768_ _2680_ _2731_ _2749_ _2750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_7_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_40_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5924__A2 _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7126__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5719_ _1034_ _1089_ _1066_ _1086_ _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
X_6699_ _2680_ _2682_ _2640_ _2683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5688__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3625__I as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5860__A1 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4663__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4456__I _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6404__A3 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7117__A1 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5391__A3 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4351__A1 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7170__C _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4050_ as2650.psl\[3\] _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_84_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4654__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xinput6 io_in[5] net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_36_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5603__A1 _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4952_ _1065_ _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3903_ _3138_ _3287_ _3438_ _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_127_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4883_ _0999_ as2650.r123_2\[2\]\[5\] _0959_ _1000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6159__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3834_ _3280_ _3369_ _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6622_ as2650.stack\[7\]\[9\] _2610_ _2611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6553_ _2490_ _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7108__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3765_ _3297_ _3300_ _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_5504_ _3228_ _1549_ _1551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6484_ _2468_ _2475_ _2489_ _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
X_3696_ _3231_ _3232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5435_ _3334_ _1484_ _1487_ _0150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_106_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6331__A2 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5366_ _1416_ _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4893__A2 _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7105_ _0308_ _0961_ _3058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_4317_ _0513_ _0514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_43_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5297_ _0413_ _1382_ _1383_ _0116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7036_ _3002_ _3004_ _3005_ _0233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4248_ _0371_ _0445_ _0439_ _0446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_28_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4179_ _0374_ _0377_ _0378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_55_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6398__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_24_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6570__A2 _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_87_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6322__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4333__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3687__A3 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6389__A2 _2395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5061__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1041 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_128_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6313__A2 _2322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4324__A1 _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5220_ _1329_ _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3758__S0 as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4875__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5151_ _0884_ _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5480__I _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6077__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4102_ _0281_ _3261_ _0302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5082_ _0522_ _1189_ _1193_ _1194_ _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_97_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5824__A1 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4627__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4033_ _3388_ _3567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_37_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5427__I1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4824__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5984_ _0695_ _1942_ _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5052__A2 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4935_ _1047_ _1048_ _1049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_36_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4866_ _0406_ _0937_ _0945_ _0984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6001__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6605_ _0701_ _2596_ _2600_ _0207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3817_ _3348_ _3352_ _3353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4797_ _3255_ _0663_ _0919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5655__I _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6536_ _2497_ _2532_ _2538_ _2539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_3748_ _3279_ _3283_ _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_107_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3679_ as2650.cycle\[3\] _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6304__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6467_ _0673_ _1558_ _1176_ _2472_ _2473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__4315__A1 _0487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5418_ as2650.r123_2\[0\]\[0\] _0912_ _1477_ _1478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA_clkbuf_leaf_45_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6398_ _2201_ _2378_ _2402_ _2405_ _2406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_47_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5349_ as2650.stack\[5\]\[11\] _1411_ _1414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_29_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7019_ _2990_ _2991_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_46_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__S0 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6435__B _2441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__I1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4734__I _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5043__A2 _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_output13_I net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6791__A2 _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3794__B _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3813__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5282__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_4_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7371__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7020__I _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6231__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5034__A2 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4720_ as2650.stack\[0\]\[6\] _0846_ _0849_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4651_ _0741_ _0798_ _0801_ _0052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5475__I as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3602_ _3137_ _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7370_ _0181_ clknet_leaf_19_wb_clk_i as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5742__B1 _1765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4582_ _0653_ _0688_ _0756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3899__A3 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6321_ as2650.stack\[2\]\[9\] _2122_ _0805_ as2650.stack\[0\]\[9\] _2331_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6252_ _0724_ _2221_ _2263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_66_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5203_ _1256_ _1262_ _1314_ _1205_ _1315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6183_ _1890_ _2194_ _2195_ _2196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_69_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5134_ _0550_ _1246_ _1247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5065_ _1055_ _1044_ _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4016_ _3482_ _3350_ _3197_ _3550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_77_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6222__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5967_ _1935_ _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6773__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4918_ _0355_ _1032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5898_ _1345_ _1911_ _1912_ _1897_ _1916_ _1917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_139_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4849_ _0929_ _0966_ _0967_ _0877_ _0968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_1_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6519_ _2458_ _3529_ _0976_ _1225_ _2522_ _2523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_107_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7244__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4729__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3633__I _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7394__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6461__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5264__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4464__I _0650_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5016__A2 _1128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4775__A1 _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5295__I _1378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6516__A2 _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3750__A2 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5255__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6870_ _1553_ _0623_ _2847_ _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_74_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5007__A2 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5821_ _1773_ _1843_ _0180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_62_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6755__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5752_ _1514_ _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4703_ _0837_ _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_30_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5683_ _0354_ _1705_ _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6507__A2 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3718__I _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7422_ _0233_ clknet_leaf_15_wb_clk_i net39 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5138__C _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4634_ _0784_ _0791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7180__A2 _3112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7267__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7353_ _0164_ clknet_leaf_12_wb_clk_i as2650.idx_ctrl\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4565_ as2650.stack\[4\]\[10\] _0737_ _0742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6304_ _1990_ _2306_ _2313_ _1966_ _2314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_144_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4496_ _0661_ _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7284_ _0095_ clknet_leaf_7_wb_clk_i as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4549__I as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6235_ _1807_ _2246_ _2247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_65_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6691__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6166_ as2650.pc\[4\] net5 _0481_ _0715_ _2179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5117_ _1225_ _1228_ _1229_ _1230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6097_ _2059_ _2061_ _2111_ _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5246__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5601__C _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5048_ _3172_ _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2806 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2817 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4284__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2828 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2839 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6999_ _2421_ _2935_ _2422_ _2972_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_0_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5954__B1 _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3980__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7171__A2 _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5182__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5182__B2 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_896 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4459__I _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6682__A1 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6674__I _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6434__A1 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6985__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4996__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6737__A2 _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4748__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_31_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3971__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7162__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5173__A1 _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5753__I _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4350_ as2650.r0\[6\] _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_141_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4369__I _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4281_ _0420_ _0477_ _0478_ _0479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_140_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6673__A1 _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6020_ _1800_ _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input4_I io_in[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6425__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6976__A2 _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5779__A3 _1804_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6922_ _2284_ _2685_ _2899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_70_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6853_ _1348_ _2674_ _2832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5804_ _3314_ _1828_ _1637_ _1829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4739__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6784_ _2763_ _0324_ _2704_ _2734_ _2735_ _2765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
X_3996_ as2650.r123\[1\]\[3\] as2650.r123_2\[1\]\[3\] _3349_ _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5735_ _1500_ _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_143_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_31_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5666_ _1702_ _0166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7153__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5164__A1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7405_ _0216_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4617_ _0749_ _0773_ _0778_ _0041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5164__B2 _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5597_ _1204_ _0657_ _1638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_85_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7336_ _0147_ clknet_leaf_1_wb_clk_i as2650.r123_2\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4548_ _0726_ _0712_ _0727_ _0023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4279__I _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7267_ _0078_ clknet_leaf_37_wb_clk_i as2650.stack\[0\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4479_ _0654_ _0657_ _0665_ _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_131_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6664__A1 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6664__B2 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6218_ _1908_ _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7198_ _0009_ clknet_leaf_1_wb_clk_i as2650.r123\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6494__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6149_ _2024_ _2161_ _2162_ _2163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5219__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6967__A2 _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_57_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2603 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2614 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2625 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2636 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_55 io_oeb[11] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2647 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_66 io_oeb[22] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2658 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_77 io_oeb[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
Xwrapped_as2650_88 io_out[33] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2669 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6719__A2 _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5059__B _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7144__A2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5155__A1 as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4902__A1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6104__B1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5458__A2 _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4917__I _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4130__A2 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6407__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6958__A2 _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4418__B1 _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7080__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5630__A2 _1491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3641__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3850_ _3385_ as2650.addr_buff\[6\] _3386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_60_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3781_ _3316_ _3241_ _3284_ _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_13_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6591__B1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5520_ _1083_ _1562_ _1563_ _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_4
XFILLER_118_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7135__A2 _3081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7184__B _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5451_ _1500_ _1502_ _1503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6894__A1 _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4402_ _0553_ _0496_ _0598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6894__B2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5382_ _1434_ _0667_ _1443_ _1444_ _1445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_114_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7121_ _3069_ _3072_ _3073_ _1572_ _3074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4333_ _0383_ _0518_ _0529_ _0530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_141_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7305__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6646__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7052_ _3002_ _3016_ _3017_ _0237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4264_ _0443_ _0457_ _0461_ _0312_ _0462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_113_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6110__A3 _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6003_ _2019_ _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4121__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4827__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4195_ _0393_ _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6949__A2 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5621__A2 _1605_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6905_ _2879_ _2881_ _2882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_54_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5658__I _3433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6836_ _2696_ _2814_ _2815_ _1691_ _0223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_24_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5909__B1 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5385__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6767_ _2638_ _2733_ _2748_ _1828_ _2749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_126_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6582__B1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3979_ _3507_ _3513_ _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_52_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5718_ _1489_ _1426_ _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6698_ _2681_ _1947_ _2682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5137__A1 _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5607__B _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5649_ _3228_ _1634_ _1687_ _1688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6885__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5688__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3699__A1 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7319_ _0130_ clknet_leaf_51_wb_clk_i as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6637__A1 _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4737__I _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output43_I net43 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A1 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4472__I _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4179__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_35_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7117__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7328__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6876__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5679__A2 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__I1 as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4351__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_69_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4647__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5851__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xinput7 io_in[6] net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyc_1
XFILLER_76_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7053__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6800__A1 _2645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7179__B _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4951_ _1064_ _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3614__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5478__I _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3902_ net10 _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4882_ _0944_ _0997_ _0998_ _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6621_ _2594_ _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_123_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3833_ _3368_ _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_119_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6552_ _2497_ _2547_ _2548_ _2553_ _2554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7108__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3764_ _3298_ _3299_ _3300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5503_ _1234_ _1547_ _1550_ _0155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3726__I _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4590__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6483_ _1172_ _2477_ _2485_ _2488_ _2489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__7345__D _0156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3695_ _3172_ _3230_ _3231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5434_ _1025_ _1477_ _1487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA_clkbuf_leaf_35_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4342__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5365_ _1426_ _1427_ _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7104_ _2465_ _3451_ _2577_ _1220_ _1785_ _3057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_87_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4316_ as2650.holding_reg\[6\] _0512_ _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_102_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5296_ _0999_ _1382_ _1383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4557__I _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7035_ net39 _3000_ _3005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4247_ _0387_ _0388_ _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_75_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6634__A4 _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5842__A2 _1267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4178_ _0294_ _0295_ _0376_ _0296_ _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_4
XFILLER_95_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5388__I _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6819_ _2665_ _2797_ _2798_ _2627_ _2799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5358__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4030__A1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3636__I _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5530__A1 net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3687__A4 _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_1211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__B1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5597__A1 _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5298__I _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__I0 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5061__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4021__A1 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6849__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4324__A2 _0520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A1 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__S1 _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5150_ _1247_ _1261_ _1262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4101_ _0297_ _0299_ _0300_ _0301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6077__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5081_ _0577_ _0585_ _0586_ _1194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5824__A2 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4032_ _3563_ _3564_ _3565_ _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_110_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6806__B _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__I0 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5588__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5983_ _1525_ _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4326__B _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4934_ _3156_ _3547_ _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5001__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_19_wb_clk_i clknet_3_3_0_wb_clk_i clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4865_ _0975_ _0897_ _0982_ _0983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6001__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6604_ as2650.stack\[7\]\[2\] _2597_ _2600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3816_ _3133_ _3350_ _3351_ _3332_ _3352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_4796_ _0917_ _0918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_118_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6535_ _1628_ _1779_ _1854_ _3537_ _2537_ _2538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3747_ _3157_ _3282_ _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_140_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6466_ _1132_ _3314_ _3230_ _2472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_134_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3678_ _3213_ _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_134_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_118_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5512__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5417_ _1476_ _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6397_ _2403_ _2404_ _2211_ _2405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5348_ _0831_ _1410_ _1413_ _0137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_82_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4079__A1 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5279_ _0858_ _1368_ _1372_ _0109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_130_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7018_ _3232_ _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3921__S1 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6170__C _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5751__A1 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4306__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4197__I _0395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_8_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5034__A3 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__B _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__B1 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4660__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4650_ as2650.stack\[2\]\[10\] _0799_ _0801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xinput10 wb_rst_i net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3601_ _3136_ _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5742__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4581_ _0754_ _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_128_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6320_ _2328_ _2329_ _2330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3899__A4 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6251_ _1773_ _2262_ _0191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_6_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5202_ _1231_ _1264_ _1265_ _1313_ _1314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_139_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6182_ _1433_ _2175_ _2195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5133_ _1203_ _1031_ _3174_ _1074_ _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_97_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5064_ _0670_ _1079_ _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3808__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7196__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4015_ _3263_ _3280_ _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6222__A2 _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5025__A3 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5966_ _0696_ _1936_ _1983_ _1691_ _0185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_52_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4917_ _0278_ _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5897_ _1896_ _1915_ _1463_ _1916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_138_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7086__C _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4848_ as2650.r0\[3\] _0935_ _0967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5733__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4779_ _3260_ _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6518_ as2650.overflow _2461_ _2521_ _1312_ _2522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_101_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6449_ _1125_ _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3914__I _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_114_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_57_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6997__B1 _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4745__I _0866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6461__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4775__A2 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5525__B _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__B1 _2961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5820_ as2650.cycle\[5\] _1842_ _1843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_90_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5751_ _3149_ _3304_ _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_97_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5486__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5963__B2 _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4702_ _0836_ _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5682_ _1715_ _1105_ _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7421_ _0232_ clknet_leaf_15_wb_clk_i net30 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_72_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4633_ _0706_ _0785_ _0790_ _0045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7352_ _0163_ clknet_leaf_21_wb_clk_i net22 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4564_ _0740_ _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6303_ _1914_ _2312_ _2313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7283_ _0094_ clknet_leaf_53_wb_clk_i as2650.ins_reg\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4495_ _0681_ _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7353__D _0164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6234_ _2243_ _2244_ _2246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6140__A1 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4297__A4 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6165_ _2177_ _2178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5116_ _3212_ _1229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6096_ _0343_ _2060_ _2111_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XTAP_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_26_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5047_ _0379_ _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_113_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4454__A1 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_34_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_2807 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2818 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2829 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6998_ _2968_ _2970_ _2701_ _2971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_129_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5949_ _0648_ _1967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_40_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4221__A4 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4233__C _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7211__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5706__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5182__A2 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7361__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6131__A1 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6176__B _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4996__A2 _1109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4748__A2 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5945__A1 _1067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3819__I _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3755__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5173__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7026__I _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4280_ _3282_ _0396_ _0403_ _0478_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_49_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6673__A2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_66_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6425__A2 _2425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6921_ _2445_ _2877_ _2898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_63_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6852_ _1272_ _0545_ _2830_ _2831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__6533__C _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5803_ _1766_ _1828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6783_ _2763_ _0324_ _2764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5936__A1 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3995_ _3472_ _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_22_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5734_ _3184_ _1636_ _1762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_17_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5665_ as2650.holding_reg\[0\] _1694_ _1701_ _1702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7384__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7404_ _0215_ clknet_leaf_34_wb_clk_i as2650.stack\[7\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4616_ as2650.stack\[3\]\[12\] _0774_ _0778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5164__A2 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5596_ _1636_ _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_129_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7335_ _0146_ clknet_leaf_64_wb_clk_i as2650.r123_2\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4547_ as2650.stack\[4\]\[7\] _0713_ _0727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7266_ _0077_ clknet_leaf_37_wb_clk_i as2650.stack\[0\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6113__A1 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4478_ _0659_ _0664_ _0665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6113__B2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6217_ _2228_ _2229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_132_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7197_ _0008_ clknet_leaf_2_wb_clk_i as2650.r123\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6148_ as2650.stack\[6\]\[5\] _1969_ _2027_ as2650.stack\[4\]\[5\] _2162_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6079_ _0709_ _2093_ _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_3327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2604 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2615 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2626 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xwrapped_as2650_56 io_oeb[12] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2637 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2648 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_67 io_oeb[23] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2659 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_78 io_oeb[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_89 io_out[34] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5927__A1 as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3639__I _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7144__A3 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6352__A1 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5155__A2 _1266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4902__A2 _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6104__A1 as2650.stack\[6\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__B2 as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4666__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_475 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7257__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A2 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6591__A1 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3780_ _3175_ _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5394__A2 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6591__B2 _2589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5450_ _3224_ _1501_ _1502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6343__A1 _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_25_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4401_ _0596_ _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6894__A2 _2652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5381_ _1081_ _1444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7120_ _1184_ _3071_ _3073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
Xclkbuf_3_2_0_wb_clk_i clknet_0_wb_clk_i clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
X_4332_ _0300_ _0524_ _0528_ _0303_ _0310_ _0529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_114_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7051_ net43 _3000_ _3017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4263_ _0458_ _0310_ _0460_ _0461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_114_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6002_ _1157_ _1430_ _2019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_80_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4194_ _0375_ _0392_ _0279_ _0393_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4121__A3 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_41_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4409__A1 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3880__A2 _3414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7071__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5082__A1 _0522_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6544__B _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4843__I _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6904_ _2670_ _2880_ _2881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_35_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_618 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6835_ net51 _2726_ _2815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5909__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_64_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5385__A2 _0656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6766_ _2739_ _2746_ _2747_ _2748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6582__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3978_ _3341_ _3414_ _3427_ _3513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_143_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6582__B2 _0989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5717_ _1744_ _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6697_ _0642_ net1 _2681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5137__A2 _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5648_ _1678_ _1682_ _1684_ _1686_ _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_136_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6885__A2 _2857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5579_ _3303_ _1014_ _1530_ _1589_ _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_117_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7318_ _0129_ clknet_leaf_51_wb_clk_i as2650.stack\[5\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7249_ _0060_ clknet_leaf_40_wb_clk_i as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4648__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6438__C _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3871__A2 _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7062__A2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output36_I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A1 _3431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4820__A1 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_10_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6325__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6876__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4887__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6628__A2 _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3832__I _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4639__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xinput8 io_in[7] net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5759__I _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5064__A1 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_17_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4950_ _3209_ _1063_ _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3614__A2 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4811__A1 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3901_ _3394_ _3431_ _3436_ _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2990 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4881_ _0467_ _0944_ _0998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6620_ _2595_ _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_60_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3832_ _3367_ _3368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6564__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6551_ _1720_ _2457_ _1583_ _2552_ _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5708__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3763_ _3185_ as2650.idx_ctrl\[0\] _3299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5502_ _1548_ _1549_ _1550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6316__A1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6482_ _2486_ _2487_ _0869_ _2488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6316__B2 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3694_ _3228_ _3229_ _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6867__A2 _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5433_ _0489_ _1484_ _1486_ _0149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_133_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4878__A1 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5364_ _0669_ _1343_ _1427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7422__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7103_ _1694_ _3055_ _1312_ _3056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4315_ _0487_ _0488_ _0491_ _0494_ _0512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_113_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5295_ _1378_ _1382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7034_ _1710_ _2996_ _3003_ _3004_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4246_ _0278_ _3420_ _0444_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_45_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4177_ _0286_ _0308_ _0376_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3853__A2 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5669__I _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5055__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A1 _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6555__A1 _2546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6818_ _1101_ _2476_ _2798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5358__A2 _0671_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6749_ _2045_ _2730_ _2731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4030__A2 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5530__A2 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_78_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3844__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5046__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__B2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5597__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4021__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7445__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6359__B _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5521__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4658__I _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4100_ _3415_ _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5080_ _0296_ _0376_ _1191_ _1192_ _1193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_97_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4031_ _3446_ _3565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_42_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5489__I as2650.addr_buff\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5037__A1 _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5588__A2 _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5982_ _1327_ _1999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_64_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4933_ _3156_ _3178_ _3422_ _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_80_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4864_ _0976_ _0895_ _0981_ _0897_ _0982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3815_ as2650.r0\[1\] _3331_ _3351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_6603_ _0841_ _2596_ _2599_ _0206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_53_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4342__B _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4795_ _0916_ _0871_ _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6534_ _1544_ _1229_ _2535_ _2536_ _1078_ _2537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6552__A4 _2553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3746_ _3281_ _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6465_ _1183_ _0920_ _1618_ _1420_ _2470_ _2471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_134_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3677_ _3144_ _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5952__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5416_ _1130_ _0925_ _1476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_134_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5512__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6396_ as2650.stack\[3\]\[11\] _1929_ _2202_ _2404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_115_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4568__I _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5347_ as2650.stack\[5\]\[10\] _1411_ _1413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_82_1035 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5278_ as2650.stack\[6\]\[11\] _1369_ _1372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4079__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7017_ _2988_ _2989_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4229_ _3345_ _0419_ _0427_ _3377_ _0428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_25_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_28_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5028__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A2 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_19_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6528__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5751__A2 _3304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5503__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6179__B _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5267__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5034__A4 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4242__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4941__I _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7029__I _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3600_ _3133_ _3135_ _3136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4580_ _0753_ _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5742__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3753__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6250_ _2219_ _1883_ _2261_ _2262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5201_ _1267_ _1311_ _1312_ _1313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_42_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4553__I0 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6181_ _2007_ _2182_ _2194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5132_ _1224_ _1230_ _1233_ _1244_ _1245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_85_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5063_ _1081_ _1175_ _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_96_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4014_ _3297_ _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_93_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6758__A1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5965_ _1885_ _1938_ _1982_ _1886_ _1983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5430__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4233__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6044__S _3325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4916_ _1029_ _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5896_ _1914_ _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_139_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4847_ _3546_ _0962_ _0964_ _0965_ _0966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6930__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5733__A2 _3305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4778_ _0358_ _0899_ _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3744__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6517_ as2650.psu\[2\] _2505_ _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3729_ _3261_ _3187_ _3262_ _3264_ _3265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_105_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7497_ net46 net17 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_49_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_31_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6448_ _2447_ _2451_ _2453_ _2454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5497__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4298__I _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6379_ _1338_ _2385_ _2386_ _2233_ _2387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3930__I _3464_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6997__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_29_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7290__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4761__I _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5078__B _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3983__A1 _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7174__A1 _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6921__A1 _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5525__C _1568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_4_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_4_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5488__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4160__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_117_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4936__I _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6988__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6988__B2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5660__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5750_ _1776_ _1647_ _1777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_76_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5963__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4701_ _0651_ _0757_ _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5681_ _1242_ _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_31_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7420_ _0231_ clknet_leaf_15_wb_clk_i net19 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4632_ as2650.stack\[2\]\[3\] _0786_ _0790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6912__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6598__I _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7351_ _0162_ clknet_leaf_21_wb_clk_i net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4563_ _0739_ _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6302_ _2308_ _2311_ _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7282_ _0093_ clknet_leaf_60_wb_clk_i as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4494_ _0675_ _0680_ _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5479__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6233_ _2243_ _2244_ _2245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4151__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6164_ as2650.pc\[6\] net7 _2177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__B1 _2253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5115_ _1226_ _1227_ _0613_ _1228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6095_ as2650.r123\[2\]\[4\] as2650.r123_2\[2\]\[4\] _3194_ _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_84_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6979__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5046_ _1149_ _3285_ _1152_ _1153_ _1158_ _1159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_100_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4067__B _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_72_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2808 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2819 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5677__I _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6997_ _1548_ _2949_ _2948_ _2969_ _2970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4581__I _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5948_ _1142_ _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5954__A2 _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7156__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5879_ _1324_ _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6903__A1 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3925__I _3459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4390__A1 as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4756__I _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3660__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_48_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6434__A3 _2440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4748__A3 _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5945__A2 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3956__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7147__A1 _1715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6920__B _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_15_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4381__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5881__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4684__A2 _0819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5633__A1 _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6920_ _1847_ _2891_ _2896_ _2516_ _2897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_94_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6851_ _2828_ _2802_ _2829_ _2830_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_62_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5802_ _0674_ _1666_ _1826_ _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA_clkbuf_leaf_54_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3994_ as2650.r0\[2\] _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6782_ _0343_ _2763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XANTENNA__5936__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5733_ _1664_ _3305_ _1761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7138__A1 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5664_ _1700_ _1701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
X_7403_ _0214_ clknet_leaf_35_wb_clk_i as2650.stack\[7\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4615_ _0745_ _0773_ _0777_ _0040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7364__D _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5595_ _3244_ _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6121__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7334_ _0145_ clknet_leaf_64_wb_clk_i as2650.r123_2\[0\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4546_ _0725_ _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4477_ _0663_ _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7265_ _0076_ clknet_leaf_44_wb_clk_i as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4124__B2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6216_ _1912_ _2222_ _2227_ _1587_ _2228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_7196_ _0007_ clknet_leaf_60_wb_clk_i as2650.r123\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XTAP_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6147_ as2650.stack\[7\]\[5\] _1968_ _1975_ as2650.stack\[5\]\[5\] _2161_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_100_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6078_ _0705_ _1986_ _2093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5029_ _0669_ _1142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_96_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2605 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2616 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2627 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2638 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_57 io_oeb[13] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2649 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_68 io_oeb[24] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_72_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xwrapped_as2650_79 io_oeb[35] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5200__I _1089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5927__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3938__A1 as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7129__A1 _0902_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3655__I as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4363__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5870__I _1888_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6104__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4115__A1 _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4666__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4486__I _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_0_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5615__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4435__B _3438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3641__A3 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6591__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_990 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4400_ _3398_ _0579_ _0593_ _0595_ _0596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4354__A1 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5380_ _1151_ _1342_ _1443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_114_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4331_ _0527_ _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5780__I _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7050_ _1728_ _2996_ _3015_ _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4262_ _0459_ _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6001_ _1240_ _0664_ _2018_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5854__A1 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4193_ _0312_ _0371_ _0382_ _0391_ _0392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_140_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5606__A1 _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5082__A2 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6903_ _1268_ _0602_ _2880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_54_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5621__A4 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6116__I _1882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7351__CLK clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6834_ _2141_ _2788_ _2809_ _2813_ _2814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_50_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5909__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5020__I _0885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6031__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6765_ _1677_ _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_50_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3977_ _3160_ _3505_ _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6582__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5716_ _1598_ _1744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4593__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6696_ _1831_ _2680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5647_ _1685_ _1499_ _1507_ _1599_ _1686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_104_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5542__B1 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5578_ _1618_ _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4896__A2 _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7317_ _0128_ clknet_leaf_50_wb_clk_i as2650.stack\[5\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4529_ _0691_ _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_104_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A1 _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7248_ _0059_ clknet_leaf_41_wb_clk_i as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A1 _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4648__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7179_ _3114_ _1704_ _1706_ _3123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_105_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A2 _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4584__A1 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6325__A2 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4336__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6696__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6089__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5533__C _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7224__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5836__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5105__I _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xinput9 io_in[8] net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__dlyb_1
XFILLER_77_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7374__CLK clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5064__A2 _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4811__A2 _0882_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3900_ _3435_ _3436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_91_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2980 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4880_ _0475_ _0946_ _0996_ _0997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2991 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3831_ _3295_ _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_92_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6380__B _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6564__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6550_ _2550_ _2551_ _1264_ _2552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3762_ as2650.idx_ctrl\[1\] _3186_ _3298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_140_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5501_ _1535_ _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6316__A2 _2316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6481_ _0913_ _3188_ _3382_ _0916_ _2487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_3693_ as2650.addr_buff\[6\] _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_12_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5432_ _1384_ _1477_ _1486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4878__A2 _0904_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5363_ _1157_ _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_138_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7102_ _1046_ _1693_ _3055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4314_ _0367_ _0510_ _0511_ _0005_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5294_ _1381_ _0115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4245_ _0383_ _0442_ _0443_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7033_ _2997_ _3461_ _3003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_132_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4176_ _0374_ _0375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_67_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6555__B _2556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5055__A2 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_3_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4802__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6004__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6817_ _0483_ _0475_ _2796_ _2797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XANTENNA__4566__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6748_ _0700_ _3543_ _2729_ _2730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6307__A2 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6679_ _3372_ _3301_ _2663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4318__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4869__A2 _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7397__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6184__C _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5046__A2 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5595__I _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6546__A2 _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4021__A3 _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4004__I net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4309__A1 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3843__I _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6359__C _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4030_ _3297_ _3471_ _3459_ _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6482__A1 _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_20_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5981_ _1989_ _1996_ _1997_ _1998_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5588__A3 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4932_ _1042_ _1045_ _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_33_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4863_ _0463_ _0889_ _0980_ _0895_ _0981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6537__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_21_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6602_ as2650.stack\[7\]\[1\] _2597_ _2599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4548__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3814_ as2650.r123\[1\]\[1\] as2650.r123_2\[1\]\[1\] _3349_ _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_4794_ _3151_ _3284_ _0916_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6533_ _2458_ _0332_ _0477_ _1225_ _3212_ _2536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3745_ _3159_ _3280_ _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6464_ _3256_ _1530_ _2469_ _2470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3676_ _3207_ _3209_ _3211_ _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_133_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5415_ _1458_ _1474_ _1475_ _0142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6170__B1 _2182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6395_ as2650.stack\[1\]\[11\] _2025_ _2027_ as2650.stack\[0\]\[11\] as2650.stack\[2\]\[11\]
+ _0754_ _2403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XANTENNA__4315__A4 _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_28_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_28_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4720__A1 as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5346_ _0827_ _1410_ _1412_ _0136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5277_ _0831_ _1368_ _1371_ _0108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_60_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6473__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7016_ _1561_ _2468_ _2984_ _2987_ _2988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
X_4228_ _3366_ _0422_ _0426_ _3371_ _0427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_29_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4159_ _0357_ _3277_ _0358_ _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_46_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6225__A1 _1652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5028__A2 _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5579__A3 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3928__I _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3762__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_11_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7282__D _0093_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5083__C _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_3_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6464__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6216__A1 _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6767__A2 _2733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4778__A1 _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6519__A2 _3529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3838__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4950__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6152__B1 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7045__I net42 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5200_ _1089_ _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_100_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6180_ _2173_ _2142_ _2193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_48_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5131_ _1234_ _1235_ _1236_ _1243_ _1244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_69_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5258__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5062_ _1032_ _1174_ _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_42_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4013_ _3170_ _3243_ _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_38_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4337__C _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_opt_2_1_wb_clk_i_I clknet_opt_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6758__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4769__A1 _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5964_ _1939_ _1981_ _1982_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4915_ _1028_ _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7367__D _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5895_ _1913_ _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3992__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4846_ _0342_ _0930_ _0962_ _0965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5194__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__B1 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4777_ _3176_ _0875_ _0899_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3744__A2 as2650.ins_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6516_ _2499_ _2515_ _2516_ _2519_ _2520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3728_ _3263_ _3242_ _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7496_ net46 net16 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4579__I _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6447_ _2452_ _3302_ _2453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3659_ _3194_ _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6694__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6378_ _1652_ _2377_ _2386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_115_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5329_ as2650.stack\[5\]\[3\] _1398_ _1402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6997__A2 _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output11_I net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3658__I _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3983__A2 _3514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4932__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4489__I _3197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4160__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6437__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6988__A2 _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_284 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4999__A1 _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5660__A2 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4952__I _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_44_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4700_ _0646_ _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3974__A2 _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5680_ _1709_ _1713_ _1714_ _0168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4631_ _0702_ _0785_ _0789_ _0044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4901__B _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7350_ _0161_ clknet_3_3_0_wb_clk_i net20 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4562_ as2650.pc\[10\] _0739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_15_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6301_ _2309_ _2310_ _2311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6125__B1 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7281_ _0092_ clknet_leaf_60_wb_clk_i as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4493_ _0678_ _3505_ _0679_ _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_144_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6676__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5479__A2 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6232_ net8 _3321_ _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_104_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__B _2807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6163_ _1888_ _2176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5114_ _3529_ _0550_ _3461_ _0976_ _1227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_97_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6094_ _1909_ _2105_ _2108_ _1104_ _2109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5045_ _1154_ _1155_ _1156_ _1157_ _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_2
XFILLER_84_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2809 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5958__I _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6996_ _2392_ _2947_ as2650.addr_buff\[4\] _2969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_129_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6600__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5947_ _1940_ _1941_ _1962_ _1964_ _1965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_0_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7156__A2 _1703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5878_ _0643_ _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_139_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_72_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4829_ _3542_ _0923_ _0949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_103_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6903__A2 _0602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_43_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_43_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4914__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1053 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4390__A2 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__A1 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6738__B _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5642__B _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6419__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5642__A2 _1529_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4772__I _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__3956__A2 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6920__C _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7147__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5817__B _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4381__A2 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4012__I _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6658__A1 _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5552__B _1584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4947__I _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3851__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5881__A2 _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7083__A1 _1234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4883__S _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6830__A1 _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5633__A2 _1672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_0_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6850_ _1100_ _0504_ _2829_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_21_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5801_ _1572_ _1825_ _1826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_90_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6781_ net29 _2761_ _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_95_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3993_ _3290_ _3526_ _3527_ _0001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5732_ _1741_ _1759_ _1760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7138__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5149__A1 _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5663_ _1696_ _1697_ _1699_ _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_7402_ _0213_ clknet_leaf_44_wb_clk_i as2650.stack\[7\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4614_ as2650.stack\[3\]\[11\] _0774_ _0777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_141_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5594_ _1563_ _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_116_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7333_ _0144_ clknet_leaf_3_wb_clk_i as2650.r123_2\[0\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4545_ _0724_ _0725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_85_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6649__A1 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7264_ _0075_ clknet_leaf_42_wb_clk_i as2650.stack\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4476_ _0660_ _0662_ _0663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_116_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7280__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__B _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6215_ _1913_ _2226_ _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4857__I as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4124__A2 _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7195_ _0006_ clknet_leaf_6_wb_clk_i as2650.r123\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__3761__I _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6146_ _1999_ _2159_ _2160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7074__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6077_ _0706_ _1984_ _2092_ _0187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_3307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6821__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5028_ _1138_ _1140_ _1141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA_input10_I wb_rst_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2606 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2617 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2628 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2639 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_58 io_oeb[14] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XFILLER_54_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xwrapped_as2650_69 io_oeb[25] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_53_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6979_ net37 _2952_ _2953_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3938__A2 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7129__A2 _1177_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3936__I _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6468__B _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4115__A2 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3671__I _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3874__A1 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5615__A2 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5598__I _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4208__S _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3641__A4 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A1 _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4007__I _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4051__A1 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_9_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4354__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A1 _1585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4330_ as2650.holding_reg\[6\] _3260_ _0526_ _0527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_5_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4261_ _0448_ _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_87_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6000_ _1239_ _2014_ _2016_ _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_119_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5854__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_input2_I io_in[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3865__A1 _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4192_ _0383_ _0386_ _0390_ _3420_ _0391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_79_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6892__I _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A2 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4409__A3 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6825__C _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6803__A1 _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6902_ _2851_ _2830_ _2878_ _2852_ _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_54_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4290__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6833_ _1915_ _2138_ _2812_ _2220_ _2813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_51_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6031__A2 _3539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6764_ _1544_ _2633_ _2745_ _2448_ _2746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3976_ _3506_ _3510_ _3511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4042__A1 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5715_ _1742_ _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4593__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6319__B1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6695_ _2659_ _2660_ _2678_ _1787_ _2679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_104_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5646_ _1519_ _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4345__A2 _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5542__A1 _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5542__B2 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5577_ _1161_ _1588_ _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_116_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7316_ _0127_ clknet_leaf_50_wb_clk_i as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4528_ _0710_ _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6288__B _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6098__A2 _2110_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4587__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7247_ _0058_ clknet_leaf_46_wb_clk_i as2650.stack\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4459_ _0645_ _0646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_120_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5845__A2 _1610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7178_ _3120_ _3121_ _3122_ _0258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_105_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7047__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6129_ _2135_ _2104_ _2143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3608__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5073__A3 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5211__I _1317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3666__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6977__I net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5533__A1 _1571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4336__A2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5814__C _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6089__A2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__A1 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7038__A1 _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6797__B1 _2762_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5121__I _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4272__A1 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2970 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__B1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2981 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2992 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4960__I _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3830_ _3365_ _3366_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4024__A1 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3761_ _3296_ _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5500_ as2650.addr_buff\[4\] _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6480_ _0896_ _0881_ _1151_ _2486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3692_ as2650.addr_buff\[5\] _3228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5431_ _0410_ _1484_ _1485_ _0148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_65_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4327__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_972 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5362_ _1418_ _1420_ _1424_ _1425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_126_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7101_ _3053_ _3054_ _1772_ _0249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_114_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4313_ as2650.r123\[2\]\[5\] _0435_ _0511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_113_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5293_ as2650.r123_2\[1\]\[4\] _0987_ _1378_ _1381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7032_ _2992_ _3002_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4244_ _0439_ _0441_ _0442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5740__B _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7199__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4175_ _0371_ _0373_ _0374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_83_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5031__I _1143_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4263__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6004__A2 _2017_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6816_ _2764_ _2794_ _2765_ _2795_ _2796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_2
XFILLER_24_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4015__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5763__A1 _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6747_ _2046_ _2699_ _2729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3959_ _3273_ _3494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6678_ _2476_ _2662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_136_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5915__B _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5629_ _1465_ _1166_ _1665_ _1427_ _1668_ _1669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4318__A2 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5515__A1 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5206__I _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4110__I _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_output41_I net41 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_30_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5506__A1 _3229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6500__I _1091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5116__I _3212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7341__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_123_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4955__I _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4493__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6234__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5980_ _1799_ _1997_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4245__A1 _0383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5588__A4 _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4931_ _1044_ _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5993__A1 _2009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_127_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5786__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4690__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4862_ _0425_ _0978_ _0888_ _0979_ _0980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_127_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_36_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6601_ _0835_ _2596_ _2598_ _0205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3813_ _3191_ _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4548__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4793_ _0914_ _0915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_140_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6532_ _3319_ _1092_ _2534_ _2535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3744_ as2650.ins_reg\[4\] as2650.ins_reg\[6\] _3162_ _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6463_ _1124_ _3285_ _2469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3675_ _3210_ _3211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_5414_ _0652_ _1457_ _1470_ _1475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6394_ _1473_ _2400_ _2401_ _2402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6170__B2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5345_ as2650.stack\[5\]\[9\] _1411_ _1412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4720__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5276_ as2650.stack\[6\]\[10\] _1369_ _1371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_29_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7015_ _3140_ _2483_ _2986_ _2987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_130_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4227_ _0425_ _3365_ _0426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6473__A2 _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4484__A1 _3138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4158_ _3244_ _3250_ _0358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_55_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6225__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4089_ _3591_ _3513_ _3579_ _3503_ _0289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_3_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5579__A4 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5696__I _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5629__C _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7214__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3944__I _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6161__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4711__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6464__A2 _1530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4475__A1 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_115_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6216__A2 _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4227__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1088 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_34_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7100__B as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A1 _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4950__A2 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6152__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6152__B2 as2650.stack\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5130_ _1237_ _1238_ _1241_ _1242_ _1243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_112_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5061_ _1173_ _1069_ _1062_ _1174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4012_ _3545_ _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_65_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6833__C _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7237__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5963_ _1743_ _1938_ _1965_ _1966_ _1980_ _1981_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5966__A1 _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4914_ _0675_ _1027_ _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_5894_ _1033_ _1325_ _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_21_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4845_ _0349_ _0883_ _0888_ _0963_ _0964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5718__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7387__CLK clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4776_ _0892_ _0889_ _0895_ _0897_ _0898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6391__B2 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6515_ _2517_ _3577_ _2518_ _2446_ _2519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3727_ as2650.ins_reg\[5\] _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_7495_ net47 net15 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3744__A3 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6143__A1 _2056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6446_ _1685_ _2452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3658_ _3193_ _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6694__A2 _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6377_ _2380_ _2384_ _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_115_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5328_ _0813_ _1397_ _1401_ _0129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5259_ _0815_ _1355_ _1360_ _0101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_75_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_21_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_17_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5420__S _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_71_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5709__A1 _1736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6382__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__B _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4932__A2 _1045_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6050__I _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6134__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6685__A2 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4696__A1 as2650.stack\[1\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6437__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4448__A1 _0434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_62_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3849__I as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3785__S _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4630_ as2650.stack\[2\]\[2\] _0786_ _0789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6373__A1 _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4561_ _0735_ _0736_ _0738_ _0025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_128_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6300_ _2266_ _2272_ _2310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7280_ _0091_ clknet_3_4_0_wb_clk_i as2650.psl\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6125__B2 _2101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4492_ _3154_ _3171_ _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6231_ _2187_ _2188_ _2242_ _2243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XANTENNA__6676__A2 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6828__C _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6162_ _2173_ _2174_ _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5113_ _0500_ _0419_ _0566_ _1226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_97_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6428__A2 _2252_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6093_ _1719_ _1893_ _1128_ as2650.addr_buff\[4\] _2107_ _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XTAP_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5044_ _3275_ _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_38_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5939__A1 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6995_ _2947_ _2967_ _2968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_53_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6061__B1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6600__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5946_ _1963_ _1948_ _1964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4611__A1 _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5877_ _0643_ _3373_ _1896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7156__A3 _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4828_ _0900_ _0948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6364__A1 _0741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4914__A2 _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4759_ _0880_ _0654_ _0881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6667__A2 _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6429_ as2650.stack\[7\]\[12\] _1929_ _0754_ as2650.stack\[6\]\[12\] _2436_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_89_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_12_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_12_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_1_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7402__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6419__A2 _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4850__A1 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3653__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_16_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5089__C _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4602__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_126_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6658__A2 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_67_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4669__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5330__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5124__I _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5094__A1 as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6830__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5800_ _1823_ _1824_ _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6780_ _2760_ _2732_ _2761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_56_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3992_ as2650.r123\[2\]\[1\] _3440_ _3527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6594__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5731_ _1321_ _1345_ _1758_ _1518_ _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_95_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6346__A1 _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5662_ _1637_ _1698_ _1097_ _1699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7401_ _0212_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4613_ _0741_ _0773_ _0776_ _0039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6897__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_650 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5593_ _1613_ _1634_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7332_ _0143_ clknet_leaf_2_wb_clk_i as2650.r123_2\[0\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_128_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4544_ as2650.pc\[7\] _0724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7425__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7263_ _0074_ clknet_leaf_40_wb_clk_i as2650.stack\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4475_ _3268_ _3217_ _0661_ _3214_ _0662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_132_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6214_ _2223_ _2225_ _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_131_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7194_ _0005_ clknet_leaf_61_wb_clk_i as2650.r123\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6145_ _2000_ _2150_ _2158_ _2159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3883__A2 _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6076_ _1985_ _2091_ _2039_ _2092_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6574__B _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5085__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6282__B1 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6821__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5027_ _0893_ _3250_ _1139_ _1140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_100_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4832__A1 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2607 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2618 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2629 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xwrapped_as2650_59 io_oeb[15] vdd vss gf180mcu_fd_sc_mcu7t5v0__tiel
XTAP_1906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_0_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6978_ _2951_ _2930_ _2952_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_0_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5929_ as2650.pc\[1\] net2 _1947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_22_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7129__A3 _3046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4348__B1 _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5560__A2 _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6468__C _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_122_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3874__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7065__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5879__I _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5615__A3 _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6576__A1 net24 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5379__A2 _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4051__A2 as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6328__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7448__CLK clknet_leaf_54_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5119__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4354__A3 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5551__A2 _1586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3862__I _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__B1 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4260_ _0447_ _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_125_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4191_ _0269_ _0389_ _0390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3865__A2 _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7056__A2 _3019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5789__I _1494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5067__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_67_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4693__I _0740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5606__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_54_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6901_ _0610_ _0602_ _2878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4290__A2 _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6832_ _2141_ _2648_ _2811_ _1428_ _2812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6567__A1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3975_ _3508_ _3509_ _3510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6763_ _2740_ _2743_ _2744_ _2745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5714_ _1439_ _1029_ _1742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6694_ _2661_ _2677_ _2678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6319__B2 as2650.stack\[4\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5790__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5645_ _1420_ _1683_ _0919_ _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_136_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5029__I _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5576_ _1527_ _1495_ _1497_ _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6569__B _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5542__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4527_ _0709_ _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7315_ _0126_ clknet_leaf_57_wb_clk_i as2650.r123\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7391__D _0202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6288__C _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6098__A3 _2112_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7246_ _0057_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4458_ _0644_ _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7177_ as2650.psu\[2\] _3120_ _1460_ _3122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4389_ _3261_ _0574_ _0585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3856__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6128_ _2141_ as2650.pc\[4\] _2104_ _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XTAP_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6059_ _1967_ _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_3127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5073__A4 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4281__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6558__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3947__I as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5230__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6479__B _2479_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3847__A2 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__B1 _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7103__B _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6797__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__B2 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_91_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4272__A2 _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6549__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2960 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__B2 _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2971 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2982 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2993 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7270__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5221__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3760_ _3295_ _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_13_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3691_ as2650.addr_buff\[7\] _3226_ _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5430_ _0999_ _1484_ _1485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_127_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3806__B _3341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4688__I _0734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5361_ _1423_ _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_58_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7100_ _3050_ _3051_ as2650.psl\[5\] _3054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4312_ _0437_ _0467_ _0509_ _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_141_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5292_ _1380_ _0114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7031_ _2989_ _2999_ _3001_ _0232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4243_ _0373_ _0385_ _0440_ _0441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6836__C _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4174_ as2650.holding_reg\[4\] _0372_ _0373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_95_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1044 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6788__A1 _1719_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4263__A2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4802__A4 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6815_ _0423_ _0399_ _2795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7386__D _0197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4015__A2 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3767__I _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5212__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6746_ _1772_ _2728_ _0220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6960__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3958_ _3488_ _3492_ _3493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6677_ _1527_ _2626_ _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3889_ _3420_ _3421_ _3424_ _3425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_109_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5982__I _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6712__A1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5628_ _1666_ _1667_ _1668_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_124_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5559_ _1598_ _1499_ _1599_ _1600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5279__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7229_ _0040_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5423__S _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5650__C _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_24_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6762__B _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5451__A1 _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4254__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_3_1_0_wb_clk_i clknet_0_wb_clk_i clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XTAP_2245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__A1 _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5203__B2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6951__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3765__A1 _3297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6703__A1 _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5506__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6937__B _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1006 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_63_wb_clk_i_I clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6656__C _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4493__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5442__A1 _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5293__I1 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4930_ _0310_ _3211_ _1043_ _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_92_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5993__A2 _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6391__C _1463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4861_ _0422_ _0977_ _0979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2790 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6600_ as2650.stack\[7\]\[0\] _2597_ _2598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_57_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3812_ _3346_ _3347_ _3348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5745__A2 _1771_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4792_ _0913_ _0871_ _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6942__A1 _2304_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6942__B2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6531_ _2533_ _2505_ _1090_ _2534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3743_ _3153_ _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3674_ _3158_ _3160_ _3210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6462_ _3433_ _1426_ _1597_ _1678_ _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_140_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5413_ _1464_ _1473_ _1474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_6393_ as2650.stack\[7\]\[11\] _0650_ _0754_ as2650.stack\[6\]\[11\] _2401_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6170__A2 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5344_ _1395_ _1411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5275_ _0827_ _1368_ _1370_ _0107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_64_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4226_ _0424_ _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7014_ _1143_ _2985_ _1620_ _1164_ _2986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6473__A3 _1086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4484__A2 _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4157_ _0356_ _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_95_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_55_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4088_ _0287_ _0288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5284__I1 _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_37_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_37_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7186__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6933__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3747__A1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6729_ _3541_ _3571_ _2712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4830__B _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5418__S _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7110__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6048__I _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5975__A2 _3462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3986__A1 _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7177__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__B1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5727__A2 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6924__B2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7189__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5127__I _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6152__A2 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_135_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3870__I _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5060_ _0336_ _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4011_ _3544_ _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5962_ _1922_ _1974_ _1978_ _1979_ _1749_ _1980_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5966__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3977__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4913_ _3170_ _3396_ _1027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7168__A1 _3114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5893_ _1034_ _1511_ _1912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4844_ _0345_ _0883_ _0963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5718__A2 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__A1 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6391__A2 _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4775_ _0896_ _3251_ _0894_ _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_119_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6514_ _2449_ _3571_ _2518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3726_ _3200_ _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_105_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7494_ net47 net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6445_ _2450_ _3391_ _2451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6143__A2 _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3657_ _3192_ _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_31_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6376_ _2381_ _2383_ _2384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5481__B _3255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5327_ as2650.stack\[5\]\[2\] _1398_ _1401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3780__I _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5258_ as2650.stack\[6\]\[3\] _1356_ _1360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5654__A1 _3185_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4209_ _3136_ _0407_ _0408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5189_ _1059_ _1284_ _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_112_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_113_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4209__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5500__I as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A1 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7159__A1 _1651_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6906__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6382__A2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4393__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4786__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5893__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5645__A1 _1420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6070__A1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_19_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6373__A2 _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5420__I1 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6241__I _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4560_ as2650.stack\[4\]\[9\] _0737_ _0738_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4491_ _0676_ _0677_ _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6125__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6230_ _1280_ _0486_ _2242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6397__B _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5884__A1 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6161_ _2141_ _2131_ _2174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_124_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5112_ _1047_ _1225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6092_ _1898_ _2100_ _2106_ _3222_ _2107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7204__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4439__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5043_ _3204_ _3212_ _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5320__I _1395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6994_ net38 _2966_ _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__5939__A2 _1956_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__B2 as2650.stack\[5\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5945_ _1067_ _1343_ _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4072__B1 _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5876_ _1890_ _1892_ _1894_ _1895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_21_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4827_ _0877_ _0947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6364__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3775__I as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4758_ _3208_ _3211_ _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_135_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_4_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3709_ as2650.ins_reg\[2\] as2650.ins_reg\[3\] _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__5990__I _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4689_ _0808_ _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_88_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6428_ as2650.stack\[5\]\[12\] _2252_ _2253_ as2650.stack\[4\]\[12\] _2435_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_88_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5875__A1 _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6100__B _2114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6359_ _2202_ _2364_ _2367_ _1749_ _2368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_103_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_27_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5627__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_52_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_124_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6052__A1 _2041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_34_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4118__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7227__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4669__A2 _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7106__B _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5341__S _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5094__A2 as2650.r0\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6291__B2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_62_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3991_ _3495_ _3525_ _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_62_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6594__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5730_ _1743_ _1748_ _1750_ _1757_ _1758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_128_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3595__I as2650.ins_reg\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5661_ _0901_ _1138_ _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_88_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6346__A2 _2354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A1 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7400_ _0211_ clknet_leaf_45_wb_clk_i as2650.stack\[7\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4612_ as2650.stack\[3\]\[10\] _0774_ _0776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4357__B2 _3547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5592_ _1627_ _1632_ _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_129_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7331_ _0142_ clknet_leaf_47_wb_clk_i as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4543_ _0722_ _0712_ _0723_ _0022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4109__A1 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7262_ _0073_ clknet_leaf_42_wb_clk_i as2650.stack\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4474_ _3180_ _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5857__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6213_ _2178_ _2181_ _2224_ _2225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_104_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7193_ _0004_ clknet_leaf_61_wb_clk_i as2650.r123\[2\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6144_ _1235_ _2151_ _2019_ _2157_ _2158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6855__B _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6075_ _2042_ _2052_ _2090_ _2037_ _2091_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XTAP_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5026_ _0305_ _3173_ _3262_ _3249_ _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_113_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7389__D _0200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2608 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2619 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6034__A1 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6977_ net36 _2951_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_80_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6585__A2 _0603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5928_ as2650.pc\[0\] net1 _1946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5859_ _1648_ _1877_ _1878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_5_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_79_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5848__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_1_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6273__A1 _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5076__A2 _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5615__A4 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5895__I _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6005__B _2021_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4339__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5000__A2 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_103_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4354__A4 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5839__A1 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5839__B2 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4190_ _0387_ _0388_ _0389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_95_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6264__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5067__A2 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6900_ net50 _2876_ _2877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_94_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_63_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6016__A1 _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6831_ _1418_ _2793_ _2810_ _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6567__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4578__A1 as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6762_ _2740_ _2743_ _2670_ _2744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3974_ _3399_ _3427_ _3413_ _3412_ _3509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
X_5713_ _1204_ _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6693_ _2668_ _2676_ _2677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6319__A2 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5644_ _0862_ _1679_ _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_15_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5575_ _1144_ _1429_ _1520_ _1555_ _1318_ _1616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7314_ _0125_ clknet_3_4_0_wb_clk_i as2650.r123\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4526_ _0708_ _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4750__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7245_ _0056_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4457_ _0643_ _0644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_131_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4089__C _3503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4502__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7176_ _1710_ _1729_ _3110_ _3121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4388_ _0578_ _0583_ _0584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_86_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6127_ _0715_ _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5058__A2 _1167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6058_ _2055_ _2063_ _2064_ _2073_ _2074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_73_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_14_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5009_ _1070_ _1119_ _1121_ _1028_ _1122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6558__A2 _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_39_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5230__A2 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6191__B1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_107_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_53_wb_clk_i_I clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_96_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3912__B _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5049__A2 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6246__B2 _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6797__A2 _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_57_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6942__C _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_17_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4272__A3 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7415__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2950 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2961 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6549__A2 _3537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2972 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2983 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2994 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5221__A2 _1331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4980__A1 _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3690_ _3182_ _3183_ _3225_ _3226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XANTENNA__5574__B _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4969__I _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6389__C _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5360_ _1422_ _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4311_ _0437_ _0508_ _0509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5291_ as2650.r123_2\[1\]\[3\] _0972_ _1378_ _1380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_114_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7030_ net30 _3000_ _3001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4242_ _0368_ _0403_ _0440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_84_1091 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4173_ _0369_ _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6237__A1 _2064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4263__A3 _0460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6814_ _1269_ _0399_ _2794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_24_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_23_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5212__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6745_ net27 _2696_ _2727_ _2728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3957_ _3491_ _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_52_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4971__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6676_ net52 _2637_ _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_108_1294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3888_ _3401_ _3406_ _3423_ _3424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5627_ _1203_ _0674_ _1667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_136_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3783__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5558_ _0862_ _1083_ _1599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_133_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4509_ as2650.pc\[1\] _0695_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
X_5489_ as2650.addr_buff\[1\] _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_133_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5279__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7228_ _0039_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_8_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_76_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7159_ _1651_ _1131_ _1072_ _1087_ _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_101_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__A1 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6228__B2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7438__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_58_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2202 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2213 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2224 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2235 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2246 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output27_I net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2257 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2268 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_41 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_15_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2279 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_70_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6400__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6951__A2 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3693__I as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7165__I _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5911__B1 _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6937__C _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_7_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_7_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6467__A1 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6219__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5690__A2 _1722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4493__A3 _0679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_64_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3868__I _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4860_ _0977_ _0978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2780 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2791 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3811_ as2650.r123\[0\]\[1\] as2650.r123\[2\]\[1\] as2650.r123_2\[0\]\[1\] as2650.r123_2\[2\]\[1\]
+ _3196_ _3323_ _3347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_60_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4791_ _3151_ _3167_ _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6942__A2 _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_53_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6530_ as2650.psu\[3\] _2533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3742_ _3276_ _3277_ _3278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_9_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6461_ _1488_ _2457_ _2464_ _2466_ _2467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6155__B1 _2168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3673_ _3208_ _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5412_ _1472_ _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6392_ as2650.stack\[5\]\[11\] _2252_ _2253_ as2650.stack\[4\]\[11\] _2400_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4181__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5343_ _1396_ _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5274_ as2650.stack\[6\]\[9\] _1369_ _1370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7024__B _2995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7013_ _3244_ _1448_ _2985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5130__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4225_ _0423_ _0424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_60_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6473__A4 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4484__A3 _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4156_ _0355_ _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6863__B _1689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_693 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4087_ _0286_ _0284_ _0287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6630__A1 _1508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3778__I _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6933__A2 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4989_ _1102_ _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3747__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6728_ _2672_ _2709_ _2710_ _2711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
XFILLER_109_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6659_ _2643_ _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6697__A1 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5942__B _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4172__A2 _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_133_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7110__A2 _3061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7260__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4475__A3 _0661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3683__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2010 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2021 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2032 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2043 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2054 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2065 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2076 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2087 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2098 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__B2 _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6924__A2 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4935__A1 _1047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_122_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6688__A1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6948__B _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5852__B _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4163__A2 _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_83_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5143__I _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_81_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6860__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4010_ _3455_ _3457_ _3544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A1 _3158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5961_ as2650.stack\[7\]\[1\] _0650_ _1921_ _1979_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_98_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3598__I as2650.ins_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_2_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4912_ _1026_ _0088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3977__A2 _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5892_ _0645_ _1889_ _1906_ _1910_ _1911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_90_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4843_ _0917_ _0962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3729__A2 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4926__A1 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4774_ _3176_ _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6513_ _1763_ _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_20_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3725_ _3260_ _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
X_7493_ net47 net13 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_140_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6679__A1 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6444_ _2449_ _2450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3656_ _3191_ _3192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7283__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6375_ _2382_ _2345_ _2383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5326_ _0841_ _1397_ _1400_ _0128_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_88_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5257_ _0813_ _1355_ _1359_ _0100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5654__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4208_ as2650.r123\[2\]\[5\] as2650.r123_2\[2\]\[5\] _3323_ _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_102_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5188_ _1295_ _1268_ _1101_ _1296_ _1299_ _1300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__3665__A1 _3195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4139_ _0336_ _0337_ _0338_ _3135_ _0339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6603__A1 _0841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3968__A2 _3354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1090 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7159__A2 _1131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4393__A2 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A1 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5228__I _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4132__I _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_0_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5893__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7095__A1 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6842__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5645__A2 _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1150 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4908__A1 _0623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4384__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4490_ _3346_ _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_143_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5333__A1 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5884__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6160_ _0720_ _2173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7086__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5111_ _1219_ _1222_ _1223_ _1224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6091_ _1337_ _2094_ _2106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XTAP_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6833__A1 _1915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5042_ _3165_ _3262_ _3250_ _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_97_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3647__A1 as2650.cycle\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6993_ net37 _2952_ _2966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_19_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6061__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5944_ _1326_ _1953_ _1961_ _1962_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_5875_ _3374_ _1893_ _1894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4826_ _0945_ _0946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4375__A2 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4757_ _3374_ _0879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5048__I _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3708_ _3243_ _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_107_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_134_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6588__B _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4688_ _0734_ _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5324__A1 _0835_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6427_ _2412_ _2433_ _2088_ _2434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3639_ _3150_ _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_108_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6358_ _2365_ _2366_ _2209_ _2367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3886__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6100__C _2020_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5309_ as2650.r123\[3\]\[3\] _1390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6289_ _2275_ _2291_ _2299_ _2300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5627__A2 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6824__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4686__I0 _0731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6052__A2 _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_21_wb_clk_i clknet_opt_1_0_wb_clk_i clknet_leaf_21_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_31_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XPHY_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_125_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__7001__A1 _2661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_13_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4366__A2 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5563__A1 _1432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6498__B _2455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_opt_2_0_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4118__A2 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7068__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5618__A2 _1160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A1 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A3 as2650.r0\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3990_ _3496_ _3524_ _3525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4054__B2 _3587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5660_ _1153_ _1657_ _1697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_90_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4611_ _0735_ _0773_ _0775_ _0038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5554__A1 _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4357__A2 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5591_ _0669_ _1249_ _1436_ _1631_ _1632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XFILLER_106_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7330_ _0141_ clknet_leaf_25_wb_clk_i as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4542_ as2650.stack\[4\]\[6\] _0713_ _0723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4109__A2 _0308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7261_ _0072_ clknet_leaf_42_wb_clk_i as2650.stack\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4473_ _3181_ _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6503__B1 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6212_ _0720_ _0557_ _2224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5857__A2 _1416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7192_ _0003_ clknet_leaf_64_wb_clk_i as2650.r123\[2\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7059__A1 _3287_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6143_ _2056_ _2156_ _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7321__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6074_ _2051_ _2074_ _2089_ _2090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_6_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_61_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6282__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5025_ _1132_ _0305_ _3396_ _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_85_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5331__I _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4293__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2609 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6034__A2 _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6976_ _1545_ _2948_ _2949_ _2950_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_54_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5927_ as2650.addr_buff\[1\] _1127_ _1422_ _1054_ _1945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__5793__A1 _3220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6990__B1 _2955_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5858_ _3271_ _1420_ _1422_ _1646_ _1877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_16_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4809_ _0914_ _0930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4348__A2 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__B1 _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5789_ _1494_ _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6111__B _2125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_43_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5848__A2 _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6273__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5241__I _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_40_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5784__A1 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6072__I _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5536__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6264__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5151__I _0884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4990__I _0357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6830_ _1102_ _2191_ _2810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_1_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_36_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4027__A1 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4578__A2 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6761_ _2711_ _2741_ _2742_ _2743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3973_ _3507_ _3508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_90_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4822__I0 _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5712_ _1739_ _1664_ _1740_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6692_ _2671_ _2673_ _2675_ _2448_ _2676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_17_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5643_ _1568_ _1259_ _1680_ _1681_ _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__6710__I _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5574_ _1323_ _1325_ _1533_ _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7313_ _0124_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4525_ as2650.pc\[4\] _0708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4750__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7244_ _0055_ clknet_leaf_48_wb_clk_i as2650.stack\[1\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_144_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4456_ _0642_ _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_137_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_132_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7175_ _1711_ _3112_ _3120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4502__A2 _0653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4387_ _0513_ _0523_ _0582_ _0583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_113_872 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6126_ _1989_ _2139_ _1997_ _2140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6057_ _2065_ _2072_ _2073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_3107 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A1 _0458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3118 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3129 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5008_ _3316_ _1120_ _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_2406 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2417 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2428 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2439 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4606__S _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4018__A1 _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_995 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7217__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6959_ _2344_ _2934_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_35_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5230__A3 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6620__I _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6191__A1 as2650.stack\[5\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5236__I _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_894 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4257__A1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4272__A4 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2940 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_75_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5839__C net9 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2951 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2962 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2973 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2984 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A1 _1436_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2995 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__B2 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_3_7_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4980__A2 _1087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6530__I as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6182__A1 _1433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5146__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4050__I as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4310_ _3310_ _0475_ _0507_ _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5290_ _1379_ _0113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4985__I _0481_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4241_ as2650.holding_reg\[5\] _0416_ _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4172_ _0368_ _0370_ _0371_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4799__A2 _3140_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_35_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6813_ net51 _2792_ _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_51_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5748__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4225__I _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6744_ _0701_ _2657_ _2725_ _2656_ _2726_ _2727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3956_ _3296_ _3445_ _3490_ _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_91_1063 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6675_ _1501_ _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3887_ _3422_ _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4971__A2 _1068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6440__I _2445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5626_ _1417_ _0657_ _1666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_137_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6173__A1 _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5557_ _0683_ _3274_ _0685_ _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__4723__A2 _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5920__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4508_ _0647_ _0692_ _0694_ _0016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5488_ _1488_ _1536_ _1539_ _0151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_117_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_132_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4439_ as2650.r123\[1\]\[1\] _0631_ _0633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_104_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7227_ _0038_ clknet_leaf_31_wb_clk_i as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4487__A1 _0669_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_59_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_104_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7158_ _1116_ _3104_ _3106_ _0254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_58_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6109_ _1921_ _2121_ _2123_ _2124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_47_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7089_ _1152_ _1178_ _3043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2203 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2214 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2225 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2236 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2247 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2258 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2269 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_42 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_14_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5739__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_30_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__4411__A1 _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6164__A1 as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5394__C _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A1 as2650.stack\[7\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5911__B2 as2650.stack\[6\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_108_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6467__A2 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4478__A1 _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6219__A2 _2142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3460 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3471 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3482 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4650__A1 as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3493 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2770 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2781 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2792 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3810_ as2650.ins_reg\[0\] _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4790_ _3431_ _0867_ _0911_ _0912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__4402__A1 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3741_ _3139_ _3205_ _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_1413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3884__I _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6460_ _2465_ _0892_ _1264_ _2466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3672_ _3162_ _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6155__A1 _1743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6155__B2 _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5411_ as2650.stack_ptr\[2\] _0648_ _1472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6391_ _1990_ _2378_ _2385_ _1915_ _1463_ _2399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XANTENNA__4705__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5342_ _1409_ _0135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_86_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7104__B1 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5273_ _1353_ _1369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4469__A1 _3215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7012_ _1566_ _1918_ _1635_ _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_4224_ net5 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_102_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5130__A2 _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4155_ _3276_ _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_68_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5969__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4086_ _0280_ _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4641__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5197__A2 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6394__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4988_ _1101_ _1102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6727_ _3463_ _3448_ _2710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3939_ _3281_ _3368_ _3474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6658_ _1455_ _3236_ _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6697__A2 net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_46_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_46_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_5609_ _0682_ _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6589_ _1254_ _2459_ _2561_ _2588_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5942__C _1145_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7405__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5514__I _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_105_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4475__A4 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4880__A1 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2000 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2011 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2022 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2033 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2044 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2055 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2066 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2077 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2088 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2099 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6385__A1 as2650.addr_buff\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5188__A2 _1268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4935__A2 _1048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6080__I _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6688__A2 _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4699__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6948__C _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7125__B _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_111_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6964__B _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_42_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6860__A2 _1418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3674__A2 _3160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6612__A2 _2603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5960_ as2650.stack\[5\]\[1\] _1975_ _1976_ as2650.stack\[4\]\[1\] as2650.stack\[6\]\[1\]
+ _1977_ _1978_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_1
XFILLER_92_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3290 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4911_ _1025_ as2650.r123_2\[2\]\[7\] _0926_ _1026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
X_5891_ _1639_ _1899_ _1907_ _1909_ _1910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_60_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4842_ _3398_ _0288_ _0311_ _0313_ _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_2
XFILLER_60_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_53_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3729__A3 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4773_ _0893_ _3285_ _0894_ _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XANTENNA__4926__A2 _1039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6512_ _1201_ _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6128__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3724_ _3259_ _3260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7492_ net46 net12 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7428__CLK clknet_leaf_2_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6679__A2 _3301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6443_ _2448_ _2449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3655_ as2650.psl\[4\] _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6374_ _2339_ _2342_ _2382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5325_ as2650.stack\[5\]\[1\] _1398_ _1400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5103__A2 _1214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5256_ as2650.stack\[6\]\[2\] _1356_ _1359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_87_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4207_ _0405_ _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5187_ as2650.psu\[2\] _3542_ _1298_ as2650.psu\[3\] _1299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5270__S _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_84_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4862__A1 _0425_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3665__A2 _3200_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4138_ as2650.r0\[4\] _3197_ _0338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XANTENNA__3789__I _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__B1 _2079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6603__A2 _2596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4069_ _0261_ _3562_ _0270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_83_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4614__A1 as2650.stack\[3\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6367__A1 _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_51_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6114__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5509__I _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4413__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6382__A4 _2389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6119__A1 as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4393__A3 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5590__A2 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_252 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_121_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7095__A2 _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4853__A1 _0961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3920__C _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6055__B1 _1815_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4605__A1 _0726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1162 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5581__A2 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_867 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5154__I _1249_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5110_ _1088_ _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7086__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6090_ _0709_ _2104_ _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5041_ _0355_ _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6833__A2 _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_112_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4844__A1 _0345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_0_wb_clk_i wb_clk_i clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_81_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6992_ _2696_ _2964_ _2965_ _0229_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_111_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5943_ _1249_ _1938_ _1954_ _1960_ _0682_ _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_34_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6349__A1 _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5874_ _0664_ _1893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_61_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7250__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4825_ _3308_ _0894_ _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4756_ _0877_ _0878_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3707_ _3159_ _3242_ _3243_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_88_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4687_ _0826_ _0063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_88_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_33_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3638_ _3173_ _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6426_ _1912_ _2415_ _2431_ _1776_ _2432_ _2433_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5324__A2 _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6357_ as2650.stack\[2\]\[10\] _1924_ _0805_ as2650.stack\[0\]\[10\] _2366_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_103_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3886__A2 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5308_ _1389_ _0121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7077__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6288_ _1818_ _2264_ _2298_ _1587_ _2299_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6285__B1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5239_ _1103_ _1339_ _1347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4835__A1 _3571_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4686__I1 as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4408__I _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_824 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4063__A2 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_38_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_73_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7001__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
Xclkbuf_leaf_61_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_61_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5938__I1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_12_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A1 _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_130_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4143__I net4 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5563__A2 _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6760__A1 _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3877__A2 _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7068__A2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_434 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5618__A3 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6815__A2 _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3629__A2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5094__A4 as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_75_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6579__A1 _2576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7273__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4054__A2 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5003__A1 _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4610_ as2650.stack\[3\]\[9\] _0774_ _0775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5590_ _0480_ _0556_ _0607_ _1630_ _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XANTENNA__5554__A2 _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4988__I _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4541_ _0721_ _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_144_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3892__I _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4472_ _0658_ _0659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6503__A1 _3283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7260_ _0071_ clknet_leaf_50_wb_clk_i as2650.stack\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6211_ as2650.pc\[7\] _0557_ _2223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_132_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5857__A3 _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7191_ _0002_ clknet_leaf_1_wb_clk_i as2650.r123\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6142_ _2154_ _2155_ _2156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7059__A2 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6806__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6708__I _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6073_ _1818_ _2042_ _2087_ _2088_ _2089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5612__I _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5024_ _1122_ _1129_ _1136_ _1137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_26_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5490__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6975_ _2392_ _2926_ _2922_ _2927_ _2949_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or4_1
XFILLER_80_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4045__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6443__I _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5926_ _3466_ _1512_ _1944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6990__A1 _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5793__A2 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4840__I1 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5857_ _0659_ _1416_ _1422_ _1876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_55_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_37_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4808_ _0900_ _0929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6742__A1 _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6742__B2 _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5788_ _1651_ _1090_ _1803_ _1814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4898__I net8 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4739_ _0860_ _0854_ _0861_ _0080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6111__C _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6409_ _2415_ _2416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7389_ _0200_ clknet_leaf_10_wb_clk_i as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_44_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5522__I _0896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7296__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5481__A1 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A1 _1336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6981__A1 _2701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5784__A2 _1803_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5536__A2 _1050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6733__A1 _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_125_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7133__B _1834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4275__A2 _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_930 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3887__I _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5224__A1 _1333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6760_ _3540_ _3566_ _3570_ _2742_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XANTENNA__6972__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3972_ _3497_ _3471_ _3507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4822__I1 as2650.r123_2\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5711_ _1568_ _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3786__A1 _3137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6691_ _1238_ _2674_ _2675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5642_ _1523_ _1529_ _0862_ _1681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5527__A2 _1564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6724__A1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5573_ _1075_ _1514_ _1436_ _1613_ _1614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XANTENNA__4511__I _0696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7312_ _0123_ clknet_leaf_55_wb_clk_i as2650.r123\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4524_ _0706_ _0692_ _0707_ _0019_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_7243_ _0054_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4455_ as2650.pc\[0\] _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4386_ _0528_ _0581_ _0582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_7174_ _2533_ _3117_ _3119_ _1798_ _0257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__4502__A3 _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__7043__B _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6125_ _2095_ _2132_ _2138_ _2101_ _1995_ _2139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XTAP_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6056_ _2066_ _2068_ _2070_ _2071_ _2072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_6_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3108 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4266__A2 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5463__A1 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3119 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5007_ _3169_ _3179_ _1120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2407 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2418 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2429 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_1706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6958_ _2626_ _2929_ _2932_ _1787_ _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6963__A1 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5909_ as2650.stack\[5\]\[0\] _0782_ _0806_ as2650.stack\[4\]\[0\] _1928_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__5230__A4 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6889_ _2861_ _2865_ _2866_ _2867_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_50_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6715__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6191__A2 _1975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4421__I as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5961__B _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7140__A1 _1056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4257__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2930 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2941 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2952 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2963 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5201__B _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2974 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6954__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2985 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5757__A2 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2996 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6706__B2 _2644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6182__A2 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4193__A1 _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3940__A1 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7131__A1 _1572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_99_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4240_ _3428_ _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5693__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4171_ _0369_ _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_132_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6237__A3 _2248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_7_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4248__A2 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_481 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5111__B _1223_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6812_ net29 _2761_ _2792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__4506__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6945__A1 net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6743_ _2622_ _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3955_ _3367_ _3489_ _3299_ _3490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_56_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4420__A2 _0604_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5765__C _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6674_ _2657_ _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3886_ _3263_ _3419_ _3422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__4971__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5625_ _1555_ _1417_ _1665_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6173__A2 _0407_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5556_ _3305_ _1504_ _1597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_3_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5920__A2 _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_464 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4507_ as2650.stack\[4\]\[0\] _0693_ _0694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7122__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5487_ _1537_ _1538_ _1539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7226_ _0037_ clknet_leaf_39_wb_clk_i as2650.stack\[3\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4438_ _3437_ _0629_ _0632_ _0008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_67_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5684__A1 _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4487__A2 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7157_ _1706_ _3103_ _3105_ _3106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_76_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4369_ _0525_ _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_98_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6108_ as2650.stack\[2\]\[4\] _2122_ _2084_ as2650.stack\[0\]\[4\] _2123_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7088_ _1444_ _1164_ _1175_ _3041_ _3042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_58_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6039_ _1715_ _1745_ _2054_ _2055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_58_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_41_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2204 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2215 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2226 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2237 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2248 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2259 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7334__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_32 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5739__A2 _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6936__A1 _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_35_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_22_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_52_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6164__A2 net7 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5911__A2 _1929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3922__A1 _3198_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7113__A1 _0445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7113__B2 _3064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6467__A3 _1176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_467 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4478__A2 _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_46_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_256 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3450 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3461 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3472 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3483 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4650__A2 _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3494 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2760 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2771 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2782 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2793 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3740_ _3274_ _3275_ _3276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_14_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5157__I net5 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3671_ _3206_ _3207_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6155__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4061__I _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5410_ _1458_ _1468_ _1471_ _0141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_6390_ _1999_ _2391_ _2397_ _2398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_127_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3913__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5341_ _0852_ as2650.stack\[5\]\[8\] _1396_ _1409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__7104__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7104__B2 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_968 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5272_ _1354_ _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7207__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A2 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7011_ net19 _2983_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5106__B _1217_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4223_ _0403_ _0421_ _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_101_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_25_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5130__A3 _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4154_ as2650.r0\[3\] _0354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7357__CLK clknet_leaf_65_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4085_ _0280_ _0284_ _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5969__A2 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6091__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_fanout51_I net31 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_102_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4236__I _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4987_ _1100_ _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6394__A2 _2400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6451__I _1263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6726_ _3463_ _3448_ _2709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3938_ as2650.ins_reg\[4\] _3264_ _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6657_ _2626_ _2636_ _2641_ _2642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3869_ _3161_ _3163_ _3405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5608_ _0683_ _0685_ _1646_ _1647_ _1648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
X_6588_ _2541_ _0597_ _2542_ _2586_ _2587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_105_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5539_ _3504_ _1580_ _1581_ _0160_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_133_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5657__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7209_ _0020_ clknet_leaf_39_wb_clk_i as2650.stack\[4\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_15_wb_clk_i clknet_3_2_0_wb_clk_i clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_47_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_8_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A1 as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2001 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_output32_I net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2012 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2023 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2034 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4632__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2045 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4146__I _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2056 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A1 _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2067 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2078 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2089 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_30_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6385__A2 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A1 _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4148__A1 _3545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1068 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4699__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6310__B _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4320__A1 _0515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6980__B _1787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3280 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4910_ _0921_ _1023_ _1024_ _1025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_3291 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5890_ _1908_ _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_33_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_55_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4841_ _0960_ _0083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2590 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4387__A1 _0513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4772_ _0875_ _0894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3729__A4 _3264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6511_ _2513_ _2514_ _2515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_1293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3723_ _3258_ _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7491_ net46 net11 vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6128__A2 as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4139__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6442_ _1500_ _2448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3654_ _3152_ _3168_ _3189_ _3190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_122_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5887__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6373_ _2339_ _1212_ _2381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_115_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_3_0_0_wb_clk_i clknet_0_wb_clk_i clknet_3_0_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_8
XFILLER_138_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5324_ _0835_ _1397_ _1399_ _0127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5639__A1 _1618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5255_ _0841_ _1355_ _1358_ _0099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_426 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4206_ _0327_ _0397_ _0398_ _3567_ _0404_ _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
X_5186_ _1297_ _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6446__I _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4137_ as2650.r123\[1\]\[4\] as2650.r123_2\[1\]\[4\] _3192_ _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_68_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4068_ _3395_ _0269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_73_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4614__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5811__A1 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_62_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5575__B1 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6709_ _1937_ _2658_ _2691_ _2692_ _2693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__6119__A2 net6 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5590__A3 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7095__A3 _3047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5260__I _1354_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6055__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6055__B2 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5802__A1 _0674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1174 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5869__A1 _1426_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5040_ _1146_ _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_100_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6991_ net37 _2624_ _1460_ _2965_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_1210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5942_ _1598_ _1958_ _1959_ _1145_ _1960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_5873_ _1891_ _1562_ _1892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_61_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4514__I as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4824_ _0866_ _0944_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4755_ _0876_ _0877_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_119_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_119_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3706_ as2650.ins_reg\[6\] as2650.ins_reg\[7\] _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4780__A1 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4686_ _0731_ as2650.stack\[1\]\[8\] _0808_ _0826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_107_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6425_ _1914_ _2425_ _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_119_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3637_ _3161_ _3173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4532__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6356_ as2650.stack\[3\]\[10\] _2206_ _0781_ as2650.stack\[1\]\[10\] _2365_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5307_ as2650.r123\[3\]\[2\] _1389_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_0_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6287_ _1029_ _2294_ _2297_ _2298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_142_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_118_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5238_ _1345_ _1329_ _1031_ _1346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_130_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5169_ as2650.psl\[5\] _0482_ _1281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6037__A1 _1084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6588__A2 _0597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4599__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5796__B1 _1821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_71_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_140_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_129_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_13_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_235 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_9_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5012__A2 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_138_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A2 _3566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_138_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_30_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_30_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_137_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5720__B1 _1746_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6276__A1 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A2 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5618__A4 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6086__I _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6028__A1 _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7418__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6579__A2 _2578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4134__S0 _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6035__B _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3801__A3 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4334__I as2650.holding_reg\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6200__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4540_ _0720_ _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_117_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_687 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4471_ as2650.addr_buff\[7\] _0658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6503__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6210_ _0724_ _2221_ _2222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7190_ _0001_ clknet_leaf_3_wb_clk_i as2650.r123\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_48_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_98_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6141_ _0481_ _0407_ _2155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6072_ _1455_ _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_135_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5023_ _1130_ _1131_ _1135_ _1136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__4509__I as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6974_ _2947_ _2393_ _2922_ _2923_ _2948_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_80_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5925_ _0695_ _1942_ _1943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5856_ _1681_ _1872_ _1874_ _1875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_142_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4807_ _0928_ _0081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5787_ _1805_ _1809_ _1810_ _1812_ _1813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_33_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4738_ as2650.stack\[0\]\[12\] _0855_ _0861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4669_ _0813_ _0809_ _0814_ _0057_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_107_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6408_ _0747_ _2414_ _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_7388_ _0199_ clknet_leaf_6_wb_clk_i as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6339_ _2176_ _2347_ _2184_ _2348_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_103_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_40_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_29_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5233__A2 _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6430__A1 _1473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4154__I as2650.r0\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A1 _3157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__B1 _0781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4744__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6497__A1 _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5713__I _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6249__A1 _2220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7240__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5869__B _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6421__A1 as2650.addr_buff\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5224__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_986 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3971_ _3404_ _3505_ _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_50_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5710_ _1738_ _0174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3786__A2 _3321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6690_ _2669_ _2674_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_31_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5641_ _1679_ _1591_ _1680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__S _1065_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1000 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5572_ _1612_ _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_7311_ _0122_ clknet_leaf_56_wb_clk_i as2650.r123\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4523_ as2650.stack\[4\]\[3\] _0693_ _0707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_129_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7242_ _0053_ clknet_leaf_38_wb_clk_i as2650.stack\[2\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4454_ _0626_ _0636_ _0641_ _0015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_1039 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7173_ _3117_ _3118_ _3119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4385_ _0531_ _3247_ _0580_ _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_131_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6124_ _2134_ _2137_ _2138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_28_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6055_ _1242_ _1513_ _1815_ as2650.addr_buff\[3\] _1210_ _2071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XTAP_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3109 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A1 _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4266__A3 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5006_ _1052_ _1118_ _1085_ _1119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_100_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5463__A2 _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2408 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2419 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6412__A1 _1649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_96_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_121_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6957_ _2639_ _2931_ _2932_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_78_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6963__A2 _2937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5908_ _1922_ _1923_ _1926_ _1927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_6888_ _1683_ _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_14_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5839_ _1578_ _1071_ _1178_ _1061_ net9 _1859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_139_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4702__I _0836_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_911 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_108_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6479__A1 _1138_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_668 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7140__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7263__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_852 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6651__A1 _2628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6651__B2 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2920 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2931 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6403__A1 _1545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2942 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2953 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2964 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2975 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2986 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2997 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A1 _3218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6706__A2 _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4717__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3940__A2 _3473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7131__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4768__B _0889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6539__I _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5443__I _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5693__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4170_ _0335_ _0339_ _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_122_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4248__A3 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3898__I _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4799__A4 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6811_ _2134_ _2790_ _2791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_63_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6945__A2 _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5748__A3 _1631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6742_ _1201_ _2719_ _2724_ _1834_ _2725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4956__A1 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3954_ _3185_ as2650.idx_ctrl\[0\] _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6673_ _1162_ _2656_ _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_3885_ _3399_ _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4522__I _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5624_ _1489_ _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5555_ _1582_ _1594_ _1596_ _0161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4506_ _0690_ _0693_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5486_ _1535_ _1538_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7122__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6449__I _1125_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5133__A1 _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7225_ _0036_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4437_ as2650.r123\[1\]\[0\] _0631_ _0632_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4397__C _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6881__A1 net32 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5684__A2 _1716_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7156_ _1333_ _1703_ _3084_ _3105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_4368_ _3444_ _0546_ _0564_ _0565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3695__A1 _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6107_ _0752_ _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7087_ _0863_ _1744_ _0303_ _3041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XTAP_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4299_ _0496_ _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6633__A1 _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6038_ _2053_ _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_73_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2205 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3998__A2 _3530_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2216 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2227 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2238 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_76_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_2249 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_77 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_42_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5528__I _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_109_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6321__B1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_49_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3440 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3451 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3462 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3473 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3484 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2750 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3495 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6927__A2 _2786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2761 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2772 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2783 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2794 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_32_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3670_ _3155_ _3206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA_clkbuf_leaf_13_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4166__A2 _3440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_63_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5340_ _0850_ _1403_ _1408_ _0134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3913__A2 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7104__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5271_ _1367_ _0106_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7010_ _2981_ _2982_ _0230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4469__A3 _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4222_ _0347_ _0317_ _0420_ _0421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5106__C _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5130__A4 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4153_ _3318_ _0332_ _0352_ _3379_ _0353_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6615__A1 _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4084_ _0281_ _0283_ _0284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_95_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5969__A3 as2650.pc\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6091__A2 _2094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4517__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_19_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6732__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_52_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4929__A1 _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4986_ _1099_ _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_51_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3937_ _3471_ _3472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6725_ _1241_ _2629_ _2627_ _2707_ _2708_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_108_1083 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6656_ _2637_ _2639_ _1828_ _1896_ _2640_ _2641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3868_ _3263_ _3404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_20_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5607_ _3149_ _3269_ _1421_ _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6587_ _2447_ _2584_ _2585_ _2586_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3799_ _3325_ _3334_ _3335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5284__S _1375_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5538_ net45 _1580_ _1470_ _1581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5106__A1 _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5469_ _3434_ _1516_ _1518_ _1520_ _1521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_121_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5657__A2 _1692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7208_ _0019_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_82_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7139_ _1071_ _1087_ _3089_ _3090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_101_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7301__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5409__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_55_wb_clk_i clknet_opt_2_1_wb_clk_i clknet_leaf_55_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__4427__I _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2002 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2013 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2024 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2035 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2046 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2057 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6909__A2 _0622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2068 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2079 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6385__A3 as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4396__A2 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7098__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A2 _1682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3950__B _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4320__A2 _0516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5721__I _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6073__A2 _2042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4084__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3270 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3281 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3292 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4840_ _0958_ as2650.r123_2\[2\]\[2\] _0959_ _0960_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XTAP_2580 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2591 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4387__A2 _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4771_ _3176_ _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5168__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6510_ _0268_ _0272_ _2514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3722_ _3257_ _3258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4139__A2 _0337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5336__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6441_ _2446_ _2447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3653_ _3177_ _3188_ _3189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6533__B1 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6372_ _0743_ _2342_ _2380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_127_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7089__A1 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5323_ as2650.stack\[5\]\[0\] _1398_ _1399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7324__CLK clknet_leaf_44_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6836__A1 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5639__A2 _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5254_ as2650.stack\[6\]\[1\] _1356_ _1358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_130_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_25_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4205_ _0402_ _0403_ _0404_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4311__A2 _0508_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5185_ net4 _1297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4136_ _3133_ _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_110_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6064__A2 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4067_ _3590_ _0267_ _3164_ _0268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4075__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_43_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5811__A2 _1153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3822__A1 _3356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__I0 _0987_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7013__A1 _3244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5575__A1 _1144_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4969_ _3359_ _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__5575__B2 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4911__S _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6708_ _2656_ _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_22_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6639_ _2623_ _2624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3889__A1 _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6827__A1 _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4866__B _0945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5541__I _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_86_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6055__A2 _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_47_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4157__I _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_572 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5566__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1186 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1197 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_106_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5716__I _1598_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4620__I _0780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5869__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6818__A1 _1101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4776__B _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_112_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_812 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6991__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6990_ _2413_ _2788_ _2955_ _2958_ _2963_ _2964_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_66_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5941_ _3465_ _1127_ _1959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_92_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5872_ as2650.addr_buff\[0\] _1891_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
Xclkbuf_leaf_0_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4823_ _0943_ _0082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5557__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4754_ _3227_ _3232_ _0875_ _0876_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3705_ _3240_ _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4780__A2 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4685_ _0726_ _0818_ _0825_ _0062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4530__I _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3636_ _3171_ _3172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6424_ _1889_ _2416_ _2419_ _2430_ _2431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_88_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6355_ _2362_ _2363_ _2364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_143_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4532__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5306_ _1388_ _0120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6286_ _2209_ _2295_ _2296_ _2297_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_66_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_959 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6285__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5237_ _1344_ _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5361__I _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4296__A1 _3193_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5168_ _1212_ _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_99_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6037__A2 _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4119_ _3298_ _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_17_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5099_ _1211_ _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5096__I0 _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5796__A1 _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_859 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5796__B2 _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6125__C _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A1 _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_33_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6760__A3 _3570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5720__A1 _1745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5720__B2 _1747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6795__C _1763_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6276__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5079__A3 _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4039__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4134__S1 _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__B2 _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_128_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6035__C _1966_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5539__A1 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6200__A2 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_128_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4350__I as2650.r0\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4470_ _3304_ _0656_ _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_128_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6140_ _2112_ _2152_ _2153_ _2154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6267__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6071_ _1030_ _2081_ _2086_ _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5022_ _1132_ _1134_ _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6019__A2 _2023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4726__S _0837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1001 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5778__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6973_ _3141_ _1617_ _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_81_645 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4525__I as2650.pc\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5924_ _0642_ _3155_ _1942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4450__A1 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5855_ _1174_ _1873_ _1032_ _1874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_139_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4806_ _0912_ as2650.r123_2\[2\]\[0\] _0927_ _0928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4202__A1 _3309_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5786_ _1811_ _1812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_119_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4737_ _0748_ _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_135_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4668_ as2650.stack\[1\]\[2\] _0810_ _0814_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6407_ _2413_ _2376_ _2414_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3619_ as2650.ins_reg\[2\] _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7387_ _0198_ clknet_3_1_0_wb_clk_i as2650.r0\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4599_ _0711_ _0766_ _0768_ _0033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_134_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6338_ _2095_ _2341_ _2346_ _2101_ _1465_ _2347_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_0_104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5091__I _1203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6269_ _2276_ _1806_ _2278_ _2280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_77_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3604__I _3139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_83_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_984 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4863__C _0895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5769__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7192__CLK clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_40_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4992__A2 _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6194__A1 as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6194__B2 as2650.stack\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5941__A1 _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4744__A2 _3272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_853 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4680__A1 _0821_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_5_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3970_ _3504_ _3208_ _3505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_90_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6185__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5640_ _1451_ _1317_ _1679_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6185__B2 _2197_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5571_ _3214_ _1497_ _1612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_79_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_106_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5932__A1 _1337_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7310_ _0121_ clknet_leaf_57_wb_clk_i as2650.r123\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4522_ _0705_ _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_129_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4453_ as2650.r123\[1\]\[7\] _0637_ _0641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7241_ _0052_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_102_1089 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7172_ _3114_ _1716_ _1717_ _3118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_125_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4384_ _3247_ _0525_ _0580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6123_ _2135_ _1270_ _2136_ _2137_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_119_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6054_ _1653_ _2049_ _2069_ _1435_ _2070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XTAP_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5005_ _1063_ _1118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_100_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6660__A2 _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5463__A3 _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_82_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2409 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6412__A2 _2230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_81_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6956_ net36 _2930_ _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4423__A1 _0618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5795__B _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5907_ _0652_ as2650.stack\[3\]\[0\] as2650.stack\[2\]\[0\] _1925_ _1926_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6887_ _2223_ _2864_ _2865_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_22_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6176__A1 _2187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5838_ _1797_ _3141_ _1798_ _1858_ _0182_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_33_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5769_ _1739_ _1082_ _1795_ _1796_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__7408__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_30_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7439_ _0250_ clknet_leaf_6_wb_clk_i as2650.carry vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_107_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_864 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6100__A1 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_461 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2910 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2921 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2932 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6403__A2 _2394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2943 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2954 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2965 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2976 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2987 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_38_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2998 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4965__A2 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A1 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_12_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5724__I _1603_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6890__A2 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4784__B _0905_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4653__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_442 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_751 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6810_ _0710_ _0425_ _2789_ _2790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_35_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_24_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_clkbuf_leaf_42_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6741_ _0700_ _2721_ _2723_ _2720_ _2724_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
X_3953_ _3442_ _3488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4956__A2 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1055 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3884_ _3419_ _3420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_91_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6672_ _1589_ _2656_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4708__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5623_ _1451_ _1517_ _1663_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_30_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5554_ _3149_ _1594_ _1595_ _1596_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_117_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4505_ _0691_ _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5485_ as2650.addr_buff\[0\] _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7122__A3 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4436_ _0630_ _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7224_ _0035_ clknet_leaf_38_wb_clk_i as2650.stack\[3\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5133__A2 _1031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7155_ as2650.psl\[1\] _3103_ _3104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5684__A3 _1717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4367_ _0548_ _0563_ _3384_ _0564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__C _2227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4892__A1 _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3695__A2 _3230_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_992 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6106_ as2650.stack\[3\]\[4\] _2075_ _2082_ as2650.stack\[1\]\[4\] _2121_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7086_ _2465_ _0604_ _2564_ _1785_ _3040_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_86_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4298_ _0495_ _0496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6094__B1 _2108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6633__A2 _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6037_ _1084_ _1423_ _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_67_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2206 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_132_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2217 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2228 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_2239 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_23 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6939_ _2308_ _2914_ _2915_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XPHY_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_23_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6149__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7230__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3758__I0 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4869__B _0986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6321__A1 as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_2_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4332__B1 _0528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6872__A2 _2848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6624__A2 _2610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3430 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_79_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3441 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3452 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3463 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3474 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3485 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__A1 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2740 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3496 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2751 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2762 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2773 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4938__A2 _1051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2784 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6324__B _2333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2795 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4623__I _0783_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_1375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_18_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5454__I _0670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_9_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5270_ _0852_ as2650.stack\[6\]\[8\] _1354_ _1367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__6312__A1 _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4221_ _3549_ _3459_ _3553_ _0306_ _0420_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_87_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4874__A1 _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4152_ _3345_ _0342_ _0351_ _3377_ _0352_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_68_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6615__A2 _2602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4083_ _0282_ _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_96_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3702__I net10 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__A1 _1338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7040__A2 _3007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7253__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4929__A2 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4985_ _0481_ _1099_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5051__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4533__I as2650.pc\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6724_ _2704_ _2705_ _2706_ _2707_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3936_ _3470_ _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1073 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6655_ _1125_ _2640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3867_ _3341_ _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_137_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5606_ _1317_ _0670_ _1341_ _1646_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6551__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6586_ _2452_ _0623_ _2585_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3798_ as2650.r123_2\[0\]\[7\] _3334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_121_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5537_ _1577_ _1578_ _1579_ _1580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_118_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6303__A1 _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5468_ _3172_ _1519_ _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_7207_ _0018_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4419_ _3450_ _0614_ _0615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_8_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4865__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5399_ _0751_ _1458_ _1461_ _1462_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7138_ _1301_ _1065_ _3089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_86_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6067__B1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6606__A2 _2597_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7069_ _3021_ _3029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_59_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4617__A1 _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5814__B1 _1827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5665__I0 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2003 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4093__A2 _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2014 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2025 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2036 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4644__S _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2047 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2058 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3840__A2 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2069 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7031__A2 _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A1 _3165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_24_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_24_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4396__A3 _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6790__A1 _1270_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5648__A3 _1684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_406 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_981 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1076 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4618__I as2650.stack_ptr\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_77_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7276__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4084__A2 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5281__A1 _0860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3260 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3271 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3282 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3293 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7022__A2 _3548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2570 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2581 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2592 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4353__I _3340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4770_ _3355_ _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5584__A2 _1615_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3721_ _3155_ _3153_ _3257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_119_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6440_ _2445_ _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3652_ _3179_ _3184_ _3187_ _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_122_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_61_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6371_ _1909_ _2375_ _2378_ _1775_ _2379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5322_ _1395_ _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__7089__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_114_222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_767 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5253_ _0835_ _1355_ _1357_ _0098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_88_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_64_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4847__A1 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4204_ _0370_ _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5184_ as2650.psu\[5\] _1296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_3_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4135_ _3346_ _0334_ _0335_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4528__I _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4066_ _3407_ _3593_ _0266_ _0267_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4075__A2 _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6743__I _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5811__A3 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3822__A2 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1094 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7013__A2 _1448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5359__I _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4968_ _3266_ _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__6772__A1 _2542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4378__A3 _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5575__A2 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6772__B2 _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6707_ _2679_ _2683_ _2690_ _1205_ _2691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4783__B1 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3919_ as2650.r0\[2\] _3196_ _3454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
X_4899_ _1013_ _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_20_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6638_ _2622_ _2623_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_137_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6524__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5327__A2 _1398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6569_ _0476_ _2555_ _2569_ _2570_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_118_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3889__A2 _3421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6827__A2 _2793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4838__A1 _0274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7299__CLK clknet_leaf_34_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_41_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4066__A2 _3593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5263__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6653__I _1617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7004__A2 _2967_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_16_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5015__A1 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1143 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1154 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4173__I _0369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1165 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A2 _1524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1198 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_8_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6515__A1 _2517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_807 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4122__B _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_6_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_83_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6818__A2 _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_106 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4829__A1 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4776__C _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_93_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_65_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_805 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4057__A2 _3445_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5254__A1 as2650.stack\[6\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5940_ _1955_ _1957_ _1958_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XFILLER_53_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_1381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3090 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5871_ _1055_ _1890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5179__I _3373_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5006__A1 _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4083__I _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4822_ _0942_ as2650.r123_2\[2\]\[1\] _0927_ _0943_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_61_573 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6754__A1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4753_ _0874_ _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_30_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3704_ _3239_ _3201_ _3240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4684_ as2650.stack\[1\]\[7\] _0819_ _0825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6423_ _1310_ _1431_ _2427_ _2429_ _2430_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_88_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3635_ _3170_ _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6354_ as2650.stack\[7\]\[10\] _2164_ _2076_ as2650.stack\[5\]\[10\] _2363_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_108_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7441__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__3740__A1 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5305_ as2650.r123\[3\]\[1\] _1388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_115_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6285_ as2650.stack\[7\]\[8\] _2206_ _2084_ as2650.stack\[4\]\[8\] _2296_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_102_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5236_ _1343_ _1344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5493__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_124_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5167_ as2650.psl\[1\] _1279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_97_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_69_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4118_ _3563_ _3536_ _0318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
X_5098_ _0557_ _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_83_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5096__I1 _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4194__S _0279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_37_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_56_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4049_ _3497_ _3445_ _3583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6993__A1 net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5796__A2 _1820_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_197 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__6745__A1 net27 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5548__A2 _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_123_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7170__A1 _1288_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5181__B1 _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5720__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_121_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_47_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4287__A2 _0480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_781 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4039__A2 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5787__A2 _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7314__CLK clknet_3_4_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6736__A1 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6736__B2 _1786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_12_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_8_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3970__A1 _3504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_3_1_wb_clk_i_I clknet_opt_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7161__A1 _1349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5462__I _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6070_ _2030_ _2083_ _2085_ _2086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_140_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_input9_I io_in[8] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5021_ _1133_ _1134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_24_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4078__I _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_26_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6972_ _2696_ _2945_ _2946_ _0228_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_19_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3710__I _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5778__A2 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6975__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6226__C _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5923_ _0695_ _0642_ _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_80_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4027__B _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5854_ _0868_ _1064_ _1873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_110_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4805_ _0926_ _0927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_107_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5785_ _1325_ _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_37_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4202__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4541__I _0721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4736_ _0858_ _0854_ _0859_ _0079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_119_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7152__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4667_ _0701_ _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6406_ as2650.pc\[11\] _2413_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3618_ _3153_ _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7386_ _0197_ clknet_leaf_0_wb_clk_i as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5702__A2 _1731_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4598_ as2650.stack\[3\]\[4\] _0767_ _0768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__3713__A1 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6337_ _2343_ _2345_ _2346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_89_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5372__I _1054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_89_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6268_ _0687_ _2278_ _2279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5219_ _1329_ _1319_ _1330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_6199_ _2202_ _2205_ _2210_ _2211_ _2212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_28_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5218__A1 _1321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7337__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3620__I _3155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5769__A2 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4441__A2 _0631_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6194__A2 _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_932 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5941__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5991__B _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7143__A1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_659 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3704__A1 _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_45_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5209__A1 _1237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6957__A1 _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_32_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4432__A2 _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_50_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5885__C _1509_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6709__A1 _1937_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6709__B2 _2692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4196__A1 _3296_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5570_ _1608_ _1609_ _1610_ _1611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5932__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4521_ _0704_ _0705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3943__A1 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7134__B2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7240_ _0051_ clknet_leaf_31_wb_clk_i as2650.stack\[2\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4452_ _0572_ _0636_ _0640_ _0014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_89_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4499__A2 _3274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7171_ _3097_ _3107_ _3117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_113_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4383_ _0578_ _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_113_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6122_ _2096_ _2099_ _2136_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_876 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_105_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6053_ _2009_ _2042_ _2069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5004_ as2650.psl\[6\] _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_54_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4671__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4536__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6948__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6955_ net35 net50 _2876_ _2930_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6412__A3 _2418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4423__A2 _0359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5620__A1 _1658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5906_ _1924_ _1925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6886_ _2178_ _2818_ _2224_ _2864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5837_ _1855_ _1590_ _1856_ _1857_ _1774_ _1858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5367__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5768_ _1774_ _1784_ _1794_ _1795_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__5923__A2 _0642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4719_ _0821_ _0845_ _0848_ _0073_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7125__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5699_ _1236_ _1578_ _1730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7438_ _0249_ clknet_leaf_60_wb_clk_i as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_135_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_102_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_49_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6198__I _1749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7369_ _0180_ clknet_leaf_17_wb_clk_i as2650.cycle\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_89_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3615__I _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_1_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__A1 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_39_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6100__A2 _2113_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4111__B2 _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5051__B _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4446__I _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2900 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6939__A1 _2308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2911 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2922 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2933 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2944 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2955 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2966 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2977 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2988 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2999 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6167__A2 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5914__A2 _1918_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_127_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5678__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_692 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4102__A1 _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_48_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A1 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A1 _1121_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4405__A2 _0600_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6740_ _2065_ _2010_ _2685_ _2722_ _2723_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3952_ _3444_ _3449_ _3486_ _3487_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_50_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4956__A3 _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6504__C _1587_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6671_ _2625_ _2653_ _2655_ _0218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_108_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3883_ _3418_ _3162_ _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_91_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5622_ _1632_ _1661_ _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_73_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_902 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5553_ _1115_ _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6520__B _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4959__C _1052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4504_ _0690_ _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5484_ _1535_ _1536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7223_ _0034_ clknet_leaf_39_wb_clk_i as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4435_ _3288_ _3327_ _3438_ _0630_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__5133__A3 _3174_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4341__A1 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7154_ _3092_ _3102_ _3103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_59_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4366_ _3318_ _0549_ _0562_ _3484_ _0563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6105_ _2024_ _2118_ _2119_ _2120_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XTAP_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7085_ _1046_ _1098_ _3038_ _3039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4297_ _0487_ _0488_ _0491_ _0494_ _0495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_80_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6094__A1 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6036_ _1989_ _2051_ _1997_ _2052_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_74_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_132_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_55_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5841__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2207 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_741 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2218 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2229 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_465 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_54_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_785 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6938_ _2309_ _2895_ _2914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XPHY_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_109_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_41_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_79 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5097__I _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6869_ _2845_ _2824_ _2846_ _2847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__3907__A1 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5825__I _1831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_135_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6321__A2 _2122_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_46_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4332__A1 _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4332__B2 _0303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A1 _1739_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3420 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_64_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3431 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3442 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3453 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3464 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3475 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2730 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2741 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3486 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6388__A2 _2377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3497 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2752 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4399__A1 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2763 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2774 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2785 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2796 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6324__C _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_144_1455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4840__S _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5735__I _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4571__A1 _0745_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_141_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6312__A2 _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4323__A1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4220_ _0418_ _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_141_267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4151_ _0345_ _3469_ _3371_ _0350_ _0351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6076__A1 _1985_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4082_ _3532_ _3534_ _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_23_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5823__A1 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4626__A2 _0786_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6379__A2 _2385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4814__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4984_ as2650.r0\[5\] _1097_ _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_23_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5051__A2 _1126_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6723_ _2704_ _2705_ _3307_ _2706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3935_ _3348_ _3352_ _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_20_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6654_ _2638_ _2639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3866_ _3399_ _3401_ _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XANTENNA__6000__A1 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_1096 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5605_ _1633_ _1644_ _1645_ _1576_ _0162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6585_ _2450_ _0603_ _2584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3797_ _3331_ _3332_ _3333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__6551__A2 _2457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_754 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5536_ _3203_ _1050_ _1579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_117_253 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_12_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_938 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5467_ _3226_ _1519_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_746 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6303__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7206_ _0017_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_132_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4418_ _0608_ _0612_ _0613_ _3452_ _0614_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_114_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5398_ _1460_ _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4865__A2 _0897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7137_ _1720_ _1567_ _3088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4349_ _0545_ _0546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1056 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7068_ _0365_ _3022_ _3028_ _0242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5665__I1 _1694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6019_ _1996_ _2023_ _2035_ _2036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_27_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2004 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2015 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2026 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2037 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2048 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2059 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6144__C _2157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5042__A2 _3262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6790__A2 _0406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_122_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
Xclkbuf_leaf_64_wb_clk_i clknet_3_0_0_wb_clk_i clknet_leaf_64_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_6_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6542__A2 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_13_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_1303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3803__I _3338_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3250 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5281__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3261 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3272 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3283 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3294 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4634__I _0784_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2560 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2571 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A1 _1280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6054__C _1435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2582 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2593 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3720_ _3255_ _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4792__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3651_ _3185_ _3186_ _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XANTENNA__5465__I _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6533__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6370_ _2377_ _2378_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_54_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5321_ _1396_ _1397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_127_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5252_ as2650.stack\[6\]\[0\] _1356_ _1357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_87_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_29_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_130_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4203_ _3565_ _0328_ _0402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5414__B _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4809__I _0914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5183_ as2650.psu\[7\] _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_68_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4134_ as2650.r123\[0\]\[4\] as2650.r123\[2\]\[4\] as2650.r123_2\[0\]\[4\] as2650.r123_2\[2\]\[4\]
+ _3331_ _0333_ _0334_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XANTENNA__7220__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4065_ _3505_ _0265_ _0266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_83_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_58_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4544__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7370__CLK clknet_leaf_19_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5024__A2 _1129_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4967_ as2650.halted _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6706_ _1937_ _2684_ _2689_ _2644_ _2690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3918_ as2650.r123\[1\]\[2\] as2650.r123_2\[1\]\[2\] _3191_ _3453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4783__A1 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4898_ net8 _1013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_6637_ _1632_ _2618_ _2621_ _2622_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
X_3849_ as2650.addr_buff\[5\] _3385_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6524__A2 _2494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6568_ _1469_ _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_4_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_98_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5519_ _1074_ _1050_ _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6499_ _1966_ _3476_ _2504_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6288__A1 _1818_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_59_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3623__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6460__A1 _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_94 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6212__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5015__A2 _1127_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1144 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_43_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1177 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5566__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__A2 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_359 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6279__A1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__B2 _1424_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7243__CLK clknet_leaf_31_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4829__A2 _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_204 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_760 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7393__CLK clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5254__A2 _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_165 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3080 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3091 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5870_ _1888_ _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6203__A1 _2175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6203__B2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4821_ _3524_ _0867_ _0941_ _0942_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XTAP_2390 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_107_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5557__A3 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4765__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4752_ _3200_ _0865_ _0874_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_144_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3703_ _3237_ _3238_ _3239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5409__B _1470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4683_ _0823_ _0818_ _0824_ _0061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5195__I _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6506__A2 _2510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6422_ _1134_ _2114_ _2428_ _2429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_135_819 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3634_ as2650.ins_reg\[4\] _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_88_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5190__A1 _1161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6353_ as2650.stack\[6\]\[10\] _1977_ _1976_ as2650.stack\[4\]\[10\] _2362_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_66_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_863 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5304_ _1387_ _0119_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_89_917 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3740__A2 _3275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6284_ as2650.stack\[6\]\[8\] _2122_ _2082_ as2650.stack\[5\]\[8\] _2295_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__4539__I as2650.pc\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5235_ _1342_ _1343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_130_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5166_ _3411_ _3372_ _0344_ _3584_ _1277_ _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_97_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_96_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4117_ _0306_ _0317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_96_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5097_ _0893_ _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4048_ _3581_ _3582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_77_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_24_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_25_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6745__A2 _2696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5999_ _1955_ _1957_ _2015_ _2016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XPHY_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_40_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3618__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_125_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7266__CLK clknet_leaf_37_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5181__B2 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5833__I _1162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6433__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6984__A2 _2957_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4184__I _3512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_16_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4995__A1 _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6736__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1066 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A1 _0336_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_63 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3970__A2 _3208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7161__A2 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_830 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA_clkbuf_leaf_61_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5020_ _0885_ _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_78_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6424__A1 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6971_ net36 _2624_ _2874_ _2946_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_93_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__A2 _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5922_ _1067_ _1326_ _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_80_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5853_ _1014_ _1523_ _1341_ _1872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__6727__A2 _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4804_ _0678_ _0925_ _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_142_1019 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5784_ _1153_ _1803_ _1810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__7289__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4735_ as2650.stack\[0\]\[11\] _0855_ _0859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4666_ _0697_ _0809_ _0812_ _0056_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6405_ _1548_ _2410_ _2411_ _2020_ _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_135_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3617_ as2650.ins_reg\[3\] _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5163__A1 _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7385_ _0196_ clknet_leaf_25_wb_clk_i as2650.pc\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4597_ _0758_ _0767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6336_ _2310_ _2307_ _2344_ _2345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__4910__A1 _0921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3713__A2 _3248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4269__I _0466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6267_ _2243_ _2244_ _2277_ _2278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XFILLER_0_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6663__A1 _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5218_ _1321_ _1322_ _1323_ _1328_ _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_131_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6198_ _1749_ _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5149_ _1257_ _1260_ _1261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6415__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5218__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_84_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4426__B1 _0599_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6966__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4977__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5828__I _1250_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_139_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3952__A2 _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6659__I _2643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_10_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_31 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4901__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6103__B1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_95_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5457__A2 _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5209__A2 _1319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6957__A2 _2931_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_91_1205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6709__A2 _2658_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4196__A2 _3470_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4520_ as2650.pc\[3\] _0704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_117_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_117_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_1047 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4451_ as2650.r123\[1\]\[6\] _0637_ _0640_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_7_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5473__I _0680_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6893__A1 _2219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4499__A3 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_660 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7170_ _1288_ _3113_ _3116_ _1691_ _0256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__6893__B2 _2870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4382_ _0575_ _0577_ _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6121_ as2650.pc\[4\] _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_115_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6052_ _2041_ _2067_ _2068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__B _2521_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5003_ _1095_ _1113_ _1114_ _1116_ _0089_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_26_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4120__A2 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5141__C _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6948__A2 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4959__A1 _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6954_ _2003_ _2925_ _2928_ _2929_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_54_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5620__A2 _1659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5905_ _0752_ _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3631__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6885_ _2701_ _2857_ _2862_ _2863_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__4552__I _0730_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5836_ _3141_ _1845_ _1857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_14_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_50_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5767_ _1785_ _1441_ _1790_ _1793_ _1794_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_108_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4718_ as2650.stack\[0\]\[5\] _0846_ _0848_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_136_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5698_ _1641_ _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7437_ _0248_ clknet_leaf_52_wb_clk_i as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4649_ _0735_ _0798_ _0800_ _0051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6884__A1 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7368_ _0179_ clknet_leaf_17_wb_clk_i as2650.cycle\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6319_ as2650.stack\[5\]\[9\] _2076_ _2079_ as2650.stack\[4\]\[9\] _2329_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_131_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7299_ _0110_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[12\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7304__CLK clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5439__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6636__A1 _1602_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1098 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_57_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2901 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2912 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2923 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2934 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2945 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2956 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2967 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2978 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2989 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4462__I _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_38_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_1260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A1 _1429_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7116__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5678__A2 _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_141_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6627__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4102__A2 _3261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_858 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5850__A2 _1163_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3861__A1 _3395_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5602__A2 _1635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3951_ _3313_ _3481_ _3485_ _3486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_63_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6073__B _2087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4372__I _0568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6670_ _2637_ _2654_ _2569_ _2655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_56_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3882_ as2650.ins_reg\[6\] _3418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_32_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5621_ _1608_ _1605_ _1656_ _1660_ _1661_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_84_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5552_ _1583_ _1564_ _1584_ _1593_ _1594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_118_936 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7107__A2 _0901_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4503_ _0651_ _0689_ _0690_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5483_ _1505_ _1508_ _1510_ _1534_ _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XFILLER_117_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7327__CLK clknet_leaf_35_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6866__A1 _2816_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4434_ _0628_ _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7222_ _0033_ clknet_leaf_39_wb_clk_i as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5133__A4 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7153_ _1333_ _1692_ _3102_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_67_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4341__A2 _0372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4365_ _3452_ _0550_ _0561_ _3479_ _0562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_113_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6104_ as2650.stack\[6\]\[4\] _2078_ _2079_ as2650.stack\[4\]\[4\] _2119_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_112_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_674 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7084_ _2561_ _1725_ _3038_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4296_ _3193_ as2650.r123\[1\]\[6\] _3326_ _0493_ _0494_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XTAP_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6094__A2 _2105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6035_ _1990_ _2042_ _2050_ _1966_ _2051_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_6_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5841__A2 _1351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3852__A1 as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2208 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2219 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7043__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_753 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1507 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1518 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_25 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1529 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_26_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6937_ _2639_ _2906_ _2912_ _1847_ _2913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XPHY_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_126_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6868_ _1213_ _0569_ _2846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5819_ _1839_ _1840_ _1842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_91_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6711__B _2694_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6799_ _1234_ _1429_ _2779_ _2780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__3907__A2 _3277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5109__A1 _1220_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_755 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6857__A1 _1832_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5046__C _1158_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_162 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6158__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_61 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4457__I _0643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5832__A2 _1675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3410 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3421 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1062 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3432 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3443 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7034__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6672__I _1589_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3454 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3465 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2720 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3476 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_60 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5045__B1 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2731 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3487 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2742 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3498 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2753 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_32_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2764 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_127_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5288__I _1374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2775 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2786 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2797 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5348__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4920__I _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4020__A1 _3549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_722 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_7 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_427 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_68_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4323__A2 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5520__A1 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4150_ _3364_ _0349_ _0350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_25_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_7_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4081_ as2650.holding_reg\[3\] _0281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__4087__A1 _0286_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5823__A2 _1823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3834__A1 _3280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_37_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6515__C _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5587__A1 _3536_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4983_ _3236_ _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5198__I _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6784__B1 _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6722_ _1239_ _3577_ _2705_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
X_3934_ _3364_ _3469_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_108_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5339__A1 as2650.stack\[5\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6653_ _1617_ _2638_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3865_ _3257_ _3295_ _3400_ _3401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6531__B _1090_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6000__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5604_ net23 _1633_ _1645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3796_ _3134_ _3332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_6584_ _2574_ _2582_ _2583_ _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5535_ _1076_ _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_106_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5466_ _1517_ _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_105_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_758 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4417_ _3584_ _3369_ _3403_ _0613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
X_7205_ _0016_ clknet_leaf_48_wb_clk_i as2650.stack\[4\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__5511__A1 _1555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4314__A2 _0510_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5397_ _1459_ _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7136_ _1772_ _3087_ _0251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_87_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4348_ _0327_ _0540_ _0542_ _3567_ _0544_ _0545_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_59_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6067__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4277__I _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7067_ as2650.r123\[0\]\[3\] _3024_ _3028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4279_ _0372_ _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_86_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5814__A2 _3268_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6018_ _1743_ _1988_ _2034_ _1919_ _2035_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_101_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3825__A1 _3359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_2005 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6492__I _2490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5610__B _1609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2016 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2027 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_54_241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2038 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2049 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_14_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1326 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1337 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1359 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_126_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4740__I _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__B _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5750__A1 _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
Xclkbuf_leaf_33_wb_clk_i clknet_3_6_0_wb_clk_i clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__5502__A1 _1548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_769 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4305__A2 _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_2_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6058__A2 _2063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5805__A2 _1825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_133_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3816__A1 _3133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7007__A1 _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3240 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7007__B2 _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4915__I _1028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3251 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_509 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3262 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3273 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3284 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3295 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5569__A1 _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2550 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2561 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2572 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2583 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6230__A2 _0486_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2594 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1860 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1871 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_144_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1882 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1893 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5584__A4 _1624_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_60_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4792__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5746__I _1595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1297 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3650_ as2650.idx_ctrl\[0\] _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XANTENNA__5741__A1 _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5320_ _1395_ _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_6_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7182__B _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6297__A2 _1211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6577__I _0574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5251_ _1353_ _1356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_47_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4202_ _3309_ _0400_ _0401_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_102_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5182_ _1288_ _1289_ _1214_ _1290_ _1293_ _1294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_123_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4133_ _3323_ _0333_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_29_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_110_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4064_ _0261_ _0262_ _0264_ _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_3_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4480__A1 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_36_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4966_ _1078_ _1079_ _1080_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_51_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6705_ _2688_ _2689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_3917_ _3344_ _3452_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4783__A2 _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4897_ _0927_ _1011_ _1012_ _0087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_137_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_22_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6636_ _1602_ _2620_ _2621_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3848_ _3383_ _3384_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5732__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6567_ _0549_ _1850_ _2559_ _2567_ _2568_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3779_ _3241_ _3314_ _3232_ _3315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_106_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5518_ _3271_ _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_133_522 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6498_ _2056_ _3524_ _2455_ _2503_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_106_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6288__A2 _2264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5449_ as2650.cycle\[6\] _1495_ _1496_ _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3904__I _3439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7119_ _0537_ _0581_ _1184_ _3071_ _3072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_130_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_12_wb_clk_i_I clknet_3_2_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5799__A1 _0655_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6436__B _1801_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7195__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6460__A2 _0892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_43_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_63_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1101 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output23_I net23 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_128_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1145 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_31_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4223__A1 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5971__A1 _1986_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_6_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5723__A1 _1489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_100_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6279__A2 _2281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_87_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_51_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_69_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6346__B _1210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_65_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7021__I _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3070 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3081 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3092 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4820_ _3492_ _0873_ _0940_ _0910_ _0941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XTAP_2380 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2391 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_18_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7177__B _1460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1690 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4751_ _0872_ _0873_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4765__A2 _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5962__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5476__I _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4380__I as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3702_ net10 _3238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4682_ as2650.stack\[1\]\[6\] _0819_ _0824_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6421_ as2650.addr_buff\[4\] _2004_ _2428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3633_ _3154_ _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_128_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5714__A1 _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6352_ _1812_ _2360_ _2361_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5190__A2 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5303_ as2650.r123\[3\]\[0\] _1387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6283_ _1921_ _2292_ _2293_ _2294_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__3724__I _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5144__C _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5234_ _1341_ _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_130_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5165_ _1254_ _1013_ _3541_ as2650.overflow _1277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_69_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_116_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4116_ _3300_ _0316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_2
XFILLER_111_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5096_ _0547_ _1208_ _1065_ _1209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_83_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4555__I as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4047_ _3579_ _3580_ _3581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XPHY_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5998_ _3462_ _1956_ _2015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_52_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4949_ _0676_ _3158_ _3504_ _1062_ _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XFILLER_123_1112 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6619_ _2608_ _0213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4508__A2 _0692_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_831 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3811__S0 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3634__I as2650.ins_reg\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_134_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6010__I _1971_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6130__A1 _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_877 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_59_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_102_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_50 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_25_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_74_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4465__I as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4444__A1 _0365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4995__A2 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_391 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_1012 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_19_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4747__A2 _0868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5944__A1 _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_30_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_7_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7210__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_1229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_143_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_1005 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_878 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_140_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4683__A1 _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6076__B _2039_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6970_ _2373_ _2658_ _2944_ _2692_ _2945_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__5632__B1 _1345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_626 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6975__A3 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1180 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5921_ _1884_ _1939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_80_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1048 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5852_ _0357_ _1869_ _1870_ _1871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_107_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4803_ _0915_ _0918_ _0921_ _0924_ _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_107_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5935__A1 _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5783_ _1639_ _1808_ _1327_ _0654_ _1809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XANTENNA__3719__I _3254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5935__B2 _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4734_ _0744_ _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_124_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4665_ as2650.stack\[1\]\[1\] _0810_ _0812_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6404_ _1542_ _1545_ _1548_ _2350_ _2411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_116_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3616_ _3151_ _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6360__A1 _2201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5163__A2 _3546_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7384_ _0195_ clknet_leaf_33_wb_clk_i as2650.pc\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4596_ _0759_ _0766_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_134_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4371__B1 _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6335_ as2650.pc\[9\] as2650.pc\[8\] _2342_ _2344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_115_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4910__A2 _1023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_115_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_748 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6266_ _0609_ _3321_ _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_103_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6765__I _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6663__A2 _1811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5217_ _0683_ _1327_ _0653_ _1328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_135_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6197_ _2207_ _2208_ _2209_ _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_85_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_40_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5148_ _0617_ _1246_ _1259_ _1260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_85_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6415__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4285__I _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5218__A3 _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5079_ _0375_ _0450_ _1189_ _1192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_72_615 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__A1 _3339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4426__B2 _3574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A2 _1074_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6179__A1 _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A1 _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_12_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7383__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6351__A1 _2054_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6351__B2 _1802_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6103__B2 as2650.stack\[5\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6675__I _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_601 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_36_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_604 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4417__A1 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_141_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_81 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_92 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4196__A3 _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6590__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5754__I _1780_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_1037 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_129_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6342__A1 _1542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4450_ _0510_ _0636_ _0639_ _0013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7174__C _1798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6893__A2 _2837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4381_ _0576_ _3338_ _0577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6120_ _2133_ _2134_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_113_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_501 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_512 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_856 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6051_ as2650.pc\[2\] _2001_ _2067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6645__A2 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_556 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__C _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_589 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5002_ _1115_ _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_85_228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_39_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7256__CLK clknet_leaf_38_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6953_ _2926_ _2922_ _2927_ _2928_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4959__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5904_ as2650.stack\[1\]\[0\] _0782_ _0806_ as2650.stack\[0\]\[0\] _1923_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_6884_ _2659_ _2860_ _2861_ _2862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5835_ _1733_ _1764_ _1847_ _1619_ _1856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_22_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5908__A1 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5766_ _1791_ _1792_ _1793_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5384__A2 _1446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4717_ _0817_ _0845_ _0847_ _0072_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5664__I _1700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5697_ _0547_ _1728_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_120_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7436_ _0247_ clknet_leaf_52_wb_clk_i as2650.ins_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4648_ as2650.stack\[2\]\[9\] _0799_ _0800_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6884__A2 _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7367_ _0178_ clknet_leaf_16_wb_clk_i as2650.cycle\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_122_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4579_ _0752_ _0753_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4895__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6318_ as2650.stack\[7\]\[9\] _2164_ _2078_ as2650.stack\[6\]\[9\] _2328_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_104_834 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_46_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_81_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7298_ _0109_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[11\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_130_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6249_ _2220_ _2258_ _2259_ _2260_ _1886_ _2261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_44_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_84_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2902 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2913 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7061__A2 _3024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2924 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2935 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_445 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2946 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5072__A1 _1183_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2957 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2968 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2979 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_13_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_1059 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5375__A2 _1431_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_775 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_786 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_458 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3689__A2 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A1 _0556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_171 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4918__I _0355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6627__A2 _2609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4638__A1 as2650.stack\[2\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6338__C _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7279__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4854__S _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3861__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3978__B _3427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7052__A2 _3016_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_21_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5063__A1 _1081_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5749__I _1511_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_264 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3950_ _3483_ _3484_ _3315_ _3485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_95_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4810__A1 _3476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6073__C _2088_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3881_ _3412_ _3414_ _3416_ _3417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_5620_ _1658_ _1659_ _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6563__A1 _1218_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5551_ _1585_ _1586_ _1592_ _1593_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5484__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_948 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4502_ _0652_ _0653_ _0688_ _0689_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XANTENNA__6315__A1 _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6315__B2 _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5482_ _1522_ _1526_ _1531_ _1533_ _1534_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_144_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7221_ _0032_ clknet_leaf_46_wb_clk_i as2650.stack\[3\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4433_ _3288_ _3327_ _0628_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4877__A1 _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7152_ _2496_ _3099_ _3101_ _0253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_99_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4341__A3 _0459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4364_ _3366_ _0556_ _0560_ _3468_ _0561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_99_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6529__B _2516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6103_ as2650.stack\[7\]\[4\] _2075_ _2076_ as2650.stack\[5\]\[4\] _2118_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_98_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_331 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4828__I _0900_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4295_ _3324_ _0492_ _0493_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7083_ _1234_ _3035_ _3037_ _0248_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_101_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A1 _0697_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6034_ _1963_ _2049_ _2050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_397 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2209 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3888__B _3423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XANTENNA__5054__A1 _3204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1508 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XTAP_1519 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6936_ _2747_ _2911_ _2912_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XPHY_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_48 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4801__A1 _3203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6867_ _1213_ _0568_ _2845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
X_5818_ _1839_ _1840_ _1841_ _0179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_52_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_50_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6554__A1 _0975_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6798_ _1417_ _2762_ _2779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_126_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5749_ _1511_ _1776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3758__I3 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6306__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7419_ _0230_ clknet_leaf_28_wb_clk_i net38 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__6857__A2 _2819_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4868__A1 _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7421__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_962 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3642__I _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_1_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4096__A2 _0265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1030 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3400 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3411 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_100_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3422 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3433 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3444 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3455 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2710 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3466 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2721 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_242 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5045__A1 _1154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2732 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3477 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5045__B2 _1157_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__B1 _1924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3488 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4473__I _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2743 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3499 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2754 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2765 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2776 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2787 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2798 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A1 _0422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5348__A2 _1410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_142_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_5_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4859__A1 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5520__A2 _1562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3921__I3 as2650.r123_2\[2\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_1_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4080_ as2650.holding_reg\[3\] _3535_ _0280_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_27_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5823__A3 _1844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3834__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4383__I _0578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4982_ _3206_ _1027_ _1096_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_63_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6721_ _2663_ _2702_ _2703_ _2704_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_2
X_3933_ _3344_ _3468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
Xclkbuf_leaf_3_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_3_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_60_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6652_ net25 _2637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3864_ as2650.holding_reg\[0\] _3245_ _3400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__6536__A1 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1065 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5603_ _1634_ _1643_ _1644_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_118_701 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6583_ _1728_ _2555_ _2569_ _2583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3795_ _3131_ _3331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__3727__I as2650.ins_reg\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5534_ _1444_ _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_756 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7444__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_12_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5465_ _1079_ _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7204_ _0015_ clknet_leaf_62_wb_clk_i as2650.r123\[1\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4416_ _0611_ _3467_ _3468_ _0612_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5511__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5396_ _3238_ _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_82_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_651 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4558__I _0691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7135_ as2650.overflow _3081_ _3086_ _3087_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4347_ _0402_ _0543_ _0544_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_101_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7066_ _0276_ _3022_ _3027_ _0241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_28_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4278_ as2650.r0\[5\] _0476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5275__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6017_ _2029_ _2033_ _2034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3825__A2 _3360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2006 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7016__A2 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2017 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2028 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5027__A1 _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2039 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1305 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1316 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6775__A1 _2625_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1327 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1338 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1349 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6919_ _2680_ _2893_ _2895_ _2896_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_74_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A1 _1685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3637__I _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_17_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5750__A2 _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_553 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA_clkbuf_leaf_41_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5502__A2 _1549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4468__I _3216_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4069__A2 _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5266__A1 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_816 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6683__I _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3816__A2 _3350_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3230 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7007__A2 _2657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3241 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3252 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4417__B _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3263 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3274 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3285 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7317__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2540 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2551 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3296 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5569__A2 _1152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2562 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2573 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2584 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1850 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2595 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1861 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_42_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_57_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4241__A2 _0416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1872 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4931__I _1044_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1883 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1894 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A1 as2650.overflow vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7019__I _2990_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6858__I _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_114_214 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5250_ _1354_ _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4201_ _0399_ _0400_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5181_ as2650.psu\[0\] _1291_ _1292_ as2650.psu\[1\] _1293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_25_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4132_ _3546_ _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_111_954 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A1 _0813_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_987 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4063_ _3258_ _0263_ _0264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_68_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_497 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5009__A1 _1070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4480__A2 _0278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_1086 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4965_ _3218_ _3147_ _1079_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_52_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6704_ _1327_ _1948_ _2685_ _2687_ _2688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_51_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_33_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6509__A1 _0438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3916_ _3369_ _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4896_ as2650.r123_2\[2\]\[6\] _0927_ _1012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3991__A1 _3495_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6635_ _1615_ _1670_ _1868_ _2619_ _2620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and4_1
XANTENNA__7182__A1 as2650.psu\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3847_ _3277_ _3382_ _3383_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_20_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_118_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6566_ _1741_ _2560_ _2566_ _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__5732__A2 _1759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3778_ _3227_ _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4997__B _1105_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5517_ _0920_ _1162_ _1560_ _1561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
X_6497_ _2499_ _2500_ _2501_ _2502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_106_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5605__C _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5448_ _3182_ _3183_ _3225_ _1500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_133_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5379_ _1440_ _1441_ _1442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_47_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7118_ as2650.holding_reg\[7\] _1160_ _3070_ _3071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_59_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7049_ _2993_ _0604_ _3015_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5799__A2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6996__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6008__I _1970_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6748__A1 _0700_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_510 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_8_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1124 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_779 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1157 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_24_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4751__I _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_54_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_790 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_840 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6920__A1 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5723__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__A1 _3266_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6678__I _2476_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_137_895 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_20 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_82 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_93 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5487__A1 _1537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_643 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_104_291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5239__A1 _1103_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__A1 _2392_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_19_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3060 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3071 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3082 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3093 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2370 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_1259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2381 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2392 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5411__A1 as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1680 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4750_ _3188_ _0871_ _0872_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_1691 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_3701_ as2650.halted _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_144_1084 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7164__A1 _1290_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4681_ _0721_ _0823_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__7164__B2 _3108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6420_ _1653_ _2425_ _2426_ _1435_ _2427_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
X_3632_ _3167_ _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6911__A1 _2885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5714__A2 _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6351_ _2054_ _2351_ _2359_ _1802_ _2360_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_127_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5492__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5190__A3 _1301_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5302_ _3328_ _1382_ _1386_ _0118_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_143_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6282_ as2650.stack\[3\]\[8\] _2206_ _2122_ as2650.stack\[2\]\[8\] _2293_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_115_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_429 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5233_ _1336_ _0680_ _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_69_610 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5164_ _0344_ _0346_ _0566_ _1272_ _1275_ _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_2
XFILLER_111_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6537__B _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4115_ _0279_ _0285_ _0314_ _0315_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_97_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5095_ _1206_ _1207_ as2650.r0\[7\] _1208_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_112_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_42_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4046_ as2650.holding_reg\[2\] _3562_ _3580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_72_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A1 _3186_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_64_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XPHY_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5997_ as2650.r123\[2\]\[2\] as2650.r123_2\[2\]\[2\] _3194_ _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_80_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5667__I _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4205__A2 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_4948_ _3159_ _3247_ _1062_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7155__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4879_ _0904_ _0994_ _0995_ _0946_ _0996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_138_648 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_53_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6618_ _0852_ as2650.stack\[7\]\[8\] _2595_ _2608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5166__B1 _0344_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5705__A2 _1734_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3716__A1 _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_134_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6549_ _1220_ _3537_ _0549_ _1223_ _2551_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XANTENNA__3915__I _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3811__S1 _3323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5469__A1 _3434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_79_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1185 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_451 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_762 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4692__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4746__I _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_102_773 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A1 _2933_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_484 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_47_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_60_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6969__B2 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7091__B1 _1179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4444__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_74_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_15_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4481__I _3279_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3955__A1 _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7146__A1 _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_607 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_139_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_629 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3707__A1 _3159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_681 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_3_3_0_wb_clk_i_I clknet_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_143_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_135_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5880__A1 _1897_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7032__I _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5632__A1 _1664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4435__A2 _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_167 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__B2 _1554_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5920_ _1937_ _0643_ _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_81_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7188__B _2496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_148 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5851_ _1442_ _1600_ _1870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4802_ _0877_ _0897_ _0922_ _0923_ _0924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_2
XANTENNA__4199__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_1119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5782_ _1807_ _1803_ _1808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5935__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4733_ _0831_ _0854_ _0857_ _0078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7137__A1 _1720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4664_ _0647_ _0809_ _0811_ _0055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5699__A1 _1236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6403_ _1545_ _2394_ _2410_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
X_3615_ _3150_ _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7383_ _0194_ clknet_leaf_33_wb_clk_i as2650.pc\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7354__D _0165_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6360__A2 _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4595_ _0706_ _0760_ _0765_ _0032_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_116_843 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6334_ _0739_ _2342_ _2343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__4371__B2 _0319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6265_ as2650.addr_buff\[0\] _2276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_88_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6112__A2 _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_857 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4123__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5216_ _1326_ _1327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6267__B _2277_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6196_ _1472_ _2209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5171__B _1278_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5147_ _1258_ _1259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_111_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_28_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_955 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5078_ _0293_ _1190_ _0288_ _3582_ _1191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_72_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__A1 _1451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_56_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_4029_ _3368_ _3354_ _3562_ _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_2
XFILLER_71_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4977__A3 _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6179__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5397__I _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_362 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5926__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_9_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__A1 _3168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6730__B _2670_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_821 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6351__A2 _2351_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_832 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_107_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_898 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_79_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6103__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4665__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5862__A1 _1660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_21 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_793 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_94_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5614__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4417__A2 _3369_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_91_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_189 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_95_1354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_885 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5100__I _1212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A1 _0537_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3756__S as2650.psl\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4196__A4 _0283_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_456 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4380_ as2650.holding_reg\[7\] _0576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_113_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_502 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_513 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_194 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_654 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6050_ _1908_ _2066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_546 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_input7_I io_in[6] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_568 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5001_ net10 _1115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4656__A2 as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5853__A1 _1014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_22_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5605__A1 _1633_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_81_402 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_947 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6952_ _2482_ _2393_ _2927_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_81_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6534__C _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5903_ _1921_ _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6883_ _1786_ _2861_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_81_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5834_ _1854_ _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_126_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5010__I _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6030__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3919__A1 as2650.r0\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5765_ _1030_ _1039_ _1778_ _1781_ _1078_ _1792_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__6550__B _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6581__A2 _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4716_ as2650.stack\[0\]\[4\] _0846_ _0847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_120_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5696_ _1700_ _1727_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7435_ _0246_ clknet_leaf_4_wb_clk_i as2650.r123\[0\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4647_ _0783_ _0799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_135_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_640 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4344__A1 _0340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7366_ _0177_ clknet_leaf_14_wb_clk_i as2650.cycle\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4578_ as2650.stack_ptr\[1\] _0751_ _0752_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_144_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4895__A2 _1001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6317_ _1812_ _2326_ _2327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_535 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7297_ _0108_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_103_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6248_ _2222_ _2260_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_130_142 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A1 _1295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6179_ _0559_ _2191_ _2020_ _2192_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_57_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6725__B _2627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_opt_3_0_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2903 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2914 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2925 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2936 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_55_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2947 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2958 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2969 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_479 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7350__CLK clknet_3_3_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6021__A1 _1988_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6021__B2 _2037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
Xclkbuf_leaf_27_wb_clk_i clknet_opt_4_0_wb_clk_i clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_90_1240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_51_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6460__B _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6572__A2 _0569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_138_220 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4583__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4335__A1 _0531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_141_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5804__B _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4886__A2 _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_684 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_71 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5835__A1 _1733_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_590 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4139__C _3135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_36_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_251 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_35_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6260__A1 _2043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5063__A2 _1175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_32_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4810__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4870__S _0959_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3880_ _3412_ _3414_ _3415_ _3416_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XANTENNA__6012__A1 _2024_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_143_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_38_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6563__A2 _0477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5550_ _1322_ _1169_ _1590_ _1591_ _1592_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_30_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4501_ _0666_ _0667_ _0674_ _0682_ _0305_ _0687_ _0688_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai33_1
XFILLER_144_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_129_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5481_ _1523_ _1532_ _3255_ _1533_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6315__A2 _2318_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7220_ _0031_ clknet_leaf_49_wb_clk_i as2650.stack\[3\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4432_ _0367_ _0626_ _0627_ _0007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_971 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_982 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7151_ _1717_ _3098_ _3100_ _3101_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
X_4363_ _0559_ _3365_ _0560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6079__A1 _0709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_310 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6102_ _1999_ _2116_ _2117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7082_ _1741_ _3035_ _3037_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4294_ as2650.r123_2\[1\]\[6\] _0492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7223__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_343 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_101_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5826__A1 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4629__A2 _0785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6033_ _2045_ _2048_ _2049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
XTAP_365 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_838 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_39_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5005__I _1063_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_27_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_6_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7373__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6251__A1 _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6264__C _1465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5054__A2 _1166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1509 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XPHY_16 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_468 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6935_ _2628_ _2908_ _2910_ _2449_ _2911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XPHY_38 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_49 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_39_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4801__A2 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6866_ _2816_ _2843_ _2844_ _0224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5817_ _1839_ _1840_ _1470_ _1841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_6797_ _1832_ _2759_ _2762_ _2639_ _2777_ _2778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XANTENNA__5675__I _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6554__A2 _2555_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4565__A1 as2650.stack\[4\]\[10\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5608__C _1647_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__S0 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5748_ _0356_ _1752_ _1631_ _1775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_2
XFILLER_124_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_124_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5679_ _0261_ _1709_ _1714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5109__A3 _0553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA_clkbuf_leaf_31_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7418_ _0229_ clknet_leaf_29_wb_clk_i net37 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7349_ _0160_ clknet_leaf_21_wb_clk_i net45 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_470 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_81_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_665 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4096__A3 _0285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3401 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_18_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3412 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3423 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3434 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2700 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3445 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_79_1146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_3456 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_17_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2711 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3467 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2722 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3478 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5045__A2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6242__A1 as2650.stack\[3\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2733 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3489 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2744 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2755 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_60_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2766 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2777 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2788 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_449 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2799 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_41_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_144_1447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_13_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6545__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_908 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_1199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7246__CLK clknet_leaf_48_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_738 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5520__A3 _1563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_974 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5808__A1 _1553_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_495 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7396__CLK clknet_leaf_49_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6481__A1 _0913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_3_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_76_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_593 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_4981_ _1058_ _1073_ _1077_ _1094_ _1095_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_51_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__6784__A2 _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3932_ _3364_ _3467_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6720_ _3463_ _3491_ _2703_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_108_1011 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_36_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6651_ _2628_ _2631_ _2635_ _2517_ _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_3863_ as2650.holding_reg\[0\] _3294_ _3246_ _3399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__5495__I _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6536__A2 _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5602_ _1121_ _1635_ _1642_ _1643_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_108_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A1 as2650.stack\[4\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6582_ _0556_ _1837_ _1855_ _0989_ _2581_ _2582_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
X_3794_ _3325_ as2650.r123\[1\]\[7\] _3327_ _3329_ _3330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XANTENNA__4332__C _0310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5533_ _1571_ _1573_ _1574_ _1576_ _0159_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_118_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_223 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5464_ _1120_ _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7203_ _0014_ clknet_leaf_6_wb_clk_i as2650.r123\[1\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4839__I _0926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4415_ _0610_ _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3743__I _3153_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5395_ _1457_ _1458_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_99_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_941 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7134_ _3082_ _3083_ _3085_ _1713_ _3081_ _3086_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_113_440 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4346_ _0495_ _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5163__C _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_685 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_836 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7065_ as2650.r123\[0\]\[2\] _3024_ _3027_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_86_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_86_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4277_ _0474_ _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_101_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6016_ _2030_ _2031_ _2032_ _2033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6472__A1 _3303_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5275__A2 _1368_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4574__I _0748_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2007 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7016__A3 _2984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2018 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A1 _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2029 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1306 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1317 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_725 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1328 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6918_ _2894_ _2895_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_23_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6527__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6849_ _1100_ _0504_ _2828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_122_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_11_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4538__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7269__CLK clknet_leaf_32_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_768 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_716 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_108_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_749 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4749__I _0870_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_40 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_2_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_51 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_123_259 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_62 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1025 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_985 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_95 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_55 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_806 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5266__A2 _1362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6463__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_24_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3220 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3231 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3242 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3253 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A1 _1913_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5018__A2 _1107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3264 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
Xclkbuf_leaf_42_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XTAP_3275 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2530 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3286 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2541 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3297 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2552 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2563 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2574 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1840 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A1 _3176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_1132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2585 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1851 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2596 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1862 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1873 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5529__B _1135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1884 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1895 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6518__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_35_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_587 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_138_1026 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__B1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4200_ _0319_ _0397_ _0398_ _3574_ _0316_ _0341_ _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi222_2
XFILLER_9_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5180_ _3464_ _1292_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_111_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4131_ _0330_ _0331_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_68_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5257__A2 _1355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_116_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4062_ _3458_ _0263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_42_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_83_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6206__A1 _0722_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4480__A3 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_64_596 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__4768__A1 _3370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4964_ _3202_ _3254_ _1078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6703_ _1944_ _2686_ _2687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__7411__CLK clknet_leaf_27_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3915_ _3317_ _3450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4895_ _0537_ _1001_ _1010_ _1011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_127_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3846_ _3227_ _3231_ _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6634_ _1526_ _1869_ _1604_ _1874_ _2619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XANTENNA__5193__A1 _1254_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6565_ _1103_ _2457_ _2563_ _2565_ _2088_ _2566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
X_3777_ _3312_ _3313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4940__A1 _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_565 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5516_ _1524_ _1558_ _1156_ _1559_ _1560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
X_6496_ _1764_ _3449_ _2501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_106_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4569__I _0744_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5174__B _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5447_ _1419_ _1498_ _1499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_105_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_248 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_99_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5378_ _1124_ _1284_ _1441_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_99_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4329_ _3259_ _0525_ _0526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7117_ _1160_ _0550_ _3070_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5248__A2 _0782_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7048_ _3012_ _2989_ _3014_ _0236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_87_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6996__A2 _2947_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_28_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_390 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6733__B _2714_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1103 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6748__A2 _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_736 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1114 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_103_75 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_35 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4759__A1 _0880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__B1 _1969_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1158 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1169 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_51_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3982__A2 _3164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_329 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_10_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5863__I _1881_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1201 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3734__A2 _3181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_524 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_3_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_88_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_771 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_622 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_281 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5239__A2 _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6987__A2 _2446_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4998__A1 _1098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3050 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3061 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3072 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_111_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3083 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6739__A2 _2698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_73_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3094 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_34_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4942__I _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2360 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2371 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2382 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2393 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_61_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5411__A2 _0648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1670 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1681 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1692 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3700_ _3152_ _3236_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_105_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_30_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4680_ _0821_ _0818_ _0822_ _0060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__7164__A2 _3109_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3631_ _3154_ _3166_ _3167_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5175__A1 _1271_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6911__A2 _2887_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6350_ _2230_ _2353_ _2355_ _2358_ _2359_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_122_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5301_ _1025_ _1375_ _1386_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_52_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_142_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6281_ as2650.stack\[1\]\[8\] _2082_ _2084_ as2650.stack\[0\]\[8\] _2292_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_5232_ _1338_ _1331_ _1340_ _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_64_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5163_ _3542_ _3546_ _1273_ _1274_ _1275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4150__A2 _0349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_964 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6427__A1 _2412_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4114_ _0311_ _0313_ _0314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_96_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_774 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5094_ as2650.r0\[6\] as2650.r0\[5\] as2650.r0\[4\] as2650.r0\[3\] _1207_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_68_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_133_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4045_ as2650.holding_reg\[2\] _3562_ _3579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XANTENNA__5013__I _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5650__A2 _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_5996_ _1893_ _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XPHY_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_80_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5402__A2 _0755_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4947_ _1060_ _1061_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_138_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_36_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3964__A2 _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_123_1125 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4878_ _0505_ _0904_ _0995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6617_ _0850_ _2602_ _2607_ _0212_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__5166__A1 _3411_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_841 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3829_ _3364_ _3365_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5166__B2 _3584_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4913__A1 _3170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3716__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6548_ _3432_ _2461_ _2549_ _1312_ _2550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_88_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7307__CLK clknet_leaf_62_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6479_ _1138_ _2478_ _2479_ _2484_ _2485_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_133_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5469__A2 _1516_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_47_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1164 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3931__I _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6969__A2 _2939_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7091__A1 _1566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7091__B2 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5641__A2 _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__3652__A1 _3179_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4762__I _3358_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1058 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_54_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5944__A3 _1961_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3955__A2 _3489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6354__B1 _2076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5593__I _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_11_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_800 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4904__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3707__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_87_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6106__B1 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_86 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A1 _2626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4002__I _3535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_888 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_65_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3841__I _3317_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_441 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5880__A2 _1898_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3891__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_66_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7082__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5632__A2 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_563 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_74_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5850_ _1517_ _1163_ _1869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__6092__C _3222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2190 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4801_ _3203_ _0880_ _0654_ _0875_ _0923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_4
XANTENNA__4199__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5781_ _1806_ _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_15_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6593__B1 _1855_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3946__A2 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4732_ as2650.stack\[0\]\[10\] _0855_ _0857_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7137__A2 _1567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5148__A1 _0617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6599__I _2594_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4663_ as2650.stack\[1\]\[0\] _0810_ _0811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_135_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3614_ _3147_ _3149_ _3150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5699__A2 _1578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6402_ _0744_ _1883_ _2408_ _2409_ _1853_ _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_116_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4594_ as2650.stack\[3\]\[3\] _0761_ _0765_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7382_ _0193_ clknet_leaf_33_wb_clk_i as2650.pc\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_6333_ _1211_ _2342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__4371__A2 _0566_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_855 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_142_140 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6264_ _1940_ _2264_ _2274_ _1465_ _2275_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_130_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_103_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5215_ _1325_ _1326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4123__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6195_ as2650.stack\[2\]\[6\] _1924_ _0805_ as2650.stack\[0\]\[6\] _2208_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_9_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5146_ _0896_ _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5171__C _1282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_474 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_69_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5077_ _3421_ _3401_ _3508_ _1190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_42_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5623__A2 _1517_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A1 _0423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4028_ _3544_ _3562_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_44_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5387__A1 _0356_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5979_ _1990_ _1988_ _1994_ _1915_ _1995_ _1996_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_2
XFILLER_55_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_139_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7128__A2 _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_958 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_424 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5139__A1 _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_21_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3926__I _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_4 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_101_1275 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_45 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_122_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4757__I _3374_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_632 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_95_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3661__I _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_121_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5862__A2 _1868_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_33 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3873__A1 _3403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__A1 _3526_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_293 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_904 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5614__A2 _1434_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_1382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_83 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5378__A1 _1124_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7119__A2 _0581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3836__I net1 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5550__A1 _1322_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_4_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_600 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_514 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_525 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4667__I _0701_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6087__C _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5000_ as2650.psu\[5\] _1095_ _1114_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_569 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5853__A2 _1523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3864__A1 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7055__A1 net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_15_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_opt_3_1_wb_clk_i clknet_opt_3_0_wb_clk_i clknet_opt_3_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_93_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A1 _2135_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6802__B2 _2720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_937 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_94_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6951_ _2885_ _2887_ _2715_ _2926_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_81_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_53_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_81_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5902_ _1920_ _1921_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6882_ _2858_ _2859_ _2860_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5369__A1 _3169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5833_ _1162_ _1854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_34_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6030__A2 net3 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3919__A2 _3196_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5764_ _1096_ _1747_ _1791_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_50_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4715_ _0836_ _0846_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6318__B1 _2078_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7365__D _0176_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3746__I _3281_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4592__A2 _0761_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5695_ _1726_ _0171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_50_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_21_wb_clk_i_I clknet_opt_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7434_ _0245_ clknet_leaf_4_wb_clk_i as2650.r123\[0\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4646_ _0784_ _0798_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_107_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4344__A2 _0321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7365_ _0176_ clknet_leaf_16_wb_clk_i as2650.cycle\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4577_ as2650.stack_ptr\[0\] _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_652 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6316_ _2054_ _2316_ _2325_ _1802_ _2326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_85_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7296_ _0107_ clknet_leaf_34_wb_clk_i as2650.stack\[6\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_118_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4577__I as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6247_ _1889_ _2229_ _1918_ _1800_ _2259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_103_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_76_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5844__A2 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6178_ _1562_ _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_57_411 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_130_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5129_ _0345_ _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_57_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2904 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3607__A1 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2915 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2926 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2937 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2948 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2959 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A1 _3282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA_clkbuf_leaf_60_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_193 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4032__A1 _3563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3656__I _3191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_254 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_788 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_438 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_107_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4335__A2 _0497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1050 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5871__I _1055_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_106_173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A2 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3846__A1 _3227_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5599__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_1190 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6207__I as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4271__A1 _0468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_90_288 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_32_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_121_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4500_ _0686_ _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5480_ _1449_ _1532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_4431_ as2650.r123\[2\]\[7\] _0435_ _0627_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4326__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5781__I _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4362_ _0558_ _0559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7150_ _1715_ _1703_ _3084_ _3100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_125_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6101_ _2000_ _2109_ _2115_ _2116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7081_ _1544_ _3035_ _3036_ _0247_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4293_ _3193_ as2650.r123\[0\]\[6\] _3333_ _0490_ _0491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_2
XFILLER_59_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_333 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_140_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5826__A2 _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6032_ _2046_ _1993_ _2047_ _2048_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XTAP_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6826__B _1677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_80_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_388 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7028__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_17 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
X_6934_ _2321_ _2909_ _2910_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5021__I _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_28 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_82_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_801 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XPHY_39 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_78_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4801__A3 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6865_ net32 _2786_ _2694_ _2844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6561__B _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_35_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4860__I _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5816_ _1568_ _1823_ _1840_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_91_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6796_ _2769_ _2776_ _2626_ _2777_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5747_ _1577_ _1774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5762__A1 _1149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3999__S1 _3349_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5678_ _1710_ _1641_ _1712_ _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_136_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7417_ _0228_ clknet_leaf_29_wb_clk_i net36 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4629_ _0697_ _0785_ _0788_ _0043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_123_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_7348_ _0159_ clknet_leaf_19_wb_clk_i net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_137_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_1_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_89_322 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_132_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7279_ _0090_ clknet_leaf_53_wb_clk_i as2650.psl\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4100__I _3415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7198__CLK clknet_leaf_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3402 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1043 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_57 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3413 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3424 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_414 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3435 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3446 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2701 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3457 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2712 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2723 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3468 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6242__A2 _0649_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3479 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_96_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2734 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2745 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2756 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_96 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2767 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2778 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2789 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5866__I _1884_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_491 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4770__I _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_14_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__B1 _1265_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_126_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5505__A1 _1235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4308__A2 _0505_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_142_706 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_116_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__5808__A2 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4945__I _0677_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5550__B _1590_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6481__A2 _3188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_23_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4492__A1 _3154_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6233__A2 _2244_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4244__A1 _0439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4980_ _1080_ _1087_ _1093_ _1094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_51_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3931_ _3465_ _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_63_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5776__I _1423_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4795__A2 _0871_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6650_ _0879_ _2634_ _2635_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_31_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_20_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3862_ _3397_ _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_5601_ net23 _1637_ _1638_ _1640_ _1641_ _1642_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_73_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4547__A2 _0713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6581_ _2491_ _2580_ _2581_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3793_ _3325_ _3328_ _3329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5532_ _1575_ _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_117_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_8_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5463_ _1513_ _1514_ _1343_ _1515_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_105_408 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7202_ _0013_ clknet_leaf_6_wb_clk_i as2650.r123\[1\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_105_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4414_ _0609_ _0610_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_126_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5394_ _1425_ _1428_ _1447_ _1456_ _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_132_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_631 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_119_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7133_ _1705_ _3084_ _1834_ _3085_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_4345_ _0541_ _0495_ _0542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__7340__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_1163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_101_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_997 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7064_ _3526_ _3022_ _3026_ _0240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_87_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4276_ _0319_ _0469_ _0472_ _0473_ _0474_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XFILLER_140_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_636 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6015_ as2650.stack\[1\]\[2\] _2025_ _1976_ as2650.stack\[0\]\[2\] _2032_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6472__A2 _0379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4483__A1 _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_55_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_100_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_27_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2008 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2019 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6224__A2 _2234_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5027__A3 _1139_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1307 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A1 _3496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1318 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_14_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1329 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_39_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6917_ _2265_ _2892_ _2894_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_70_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5686__I _1289_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1123 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6848_ _2662_ _2825_ _2826_ _2667_ _2827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_10_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4538__A2 _0712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6779_ net28 _2760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_109_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_213 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_920 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_791 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_30 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_46_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_942 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_12 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4710__A2 _0839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_174 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_848 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_77_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_967 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6463__A2 _3285_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_86_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3210 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_20_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_3221 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3232 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3243 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3254 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6215__A2 _2226_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3265 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2520 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3276 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2531 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2542 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3287 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3298 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_33_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2553 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2564 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A1 _0699_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1830 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4777__A2 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2575 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5596__I _1636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1841 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2586 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_60_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1852 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2597 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1863 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_18_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_13_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1874 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1885 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1245 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1896 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7213__CLK clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5726__A1 _1258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_31_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5741__A4 _1768_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7363__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6151__A1 as2650.stack\[3\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_750 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_69_826 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_123_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4130_ _3389_ _0317_ _0318_ _0327_ _0329_ _0330_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_4
XFILLER_68_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_934 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_271 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4675__I _0807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4061_ _3257_ _0262_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_37_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_114_1082 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6206__A2 _1936_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_873 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4963_ _0868_ _1074_ _1076_ _1063_ _1077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XANTENNA__4768__A2 _0886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5965__A1 _1885_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6702_ _1807_ _2660_ _2686_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_36_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3914_ _3448_ _3449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_4894_ _1001_ _1008_ _1009_ _1010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_138_809 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6633_ _2616_ _2617_ _1067_ _1326_ _2618_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_3845_ _3311_ _3313_ _3315_ _3380_ _3381_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6914__B1 _2890_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6564_ _2465_ _0604_ _2564_ _1232_ _2565_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5193__A2 _0611_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3776_ _3251_ _3278_ _3312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5515_ _1051_ _1120_ _1559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_121_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4940__A2 _3219_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6495_ _1685_ _3492_ _2500_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_105_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5446_ _3224_ _1495_ _1497_ _1498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_47_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5377_ _1027_ _1038_ _1440_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_102_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7116_ _0536_ _0581_ _3066_ _3067_ _3068_ _3069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_99_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4328_ _0512_ _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6445__A2 _3391_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4585__I _0758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7047_ _0476_ _2991_ _2988_ _3013_ _3014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_4259_ _0444_ _0453_ _0456_ _0457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and3_1
XFILLER_101_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_477 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6733__C _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1115 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7236__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1137 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4759__A2 _0654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_58 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5956__B2 as2650.stack\[2\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_42_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1148 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_19_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_93_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A1 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7386__CLK clknet_leaf_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6381__A1 as2650.addr_buff\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_1104 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3734__A3 _3269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3664__I _3199_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7283__D _0094_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_897 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6040__I _1453_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6133__A1 _1653_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_536 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_84 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_2_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A1 _0831_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_105_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_26_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_61_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_72 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4495__I _0681_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_120_764 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_77_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_24_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_19_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_114 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3040 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_1353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3051 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_37_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_4_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_92_169 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3062 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_361 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3073 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3084 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3095 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2350 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2361 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A1 _1940_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_2_1092 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2372 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2383 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2394 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1660 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1671 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1682 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4163__C _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1693 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_144_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_820 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3630_ _3157_ _3158_ _3165_ _3166_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XANTENNA__6372__A1 _0743_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5175__A2 _1276_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_341 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__4922__A2 _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5300_ _0492_ _1382_ _1385_ _0117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_66_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6280_ _2064_ _2290_ _2291_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_45_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5231_ _1241_ _1339_ _1340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_103_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_9_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5162_ _0677_ _0269_ _1068_ _1106_ _1274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand4_1
XFILLER_111_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4113_ _0312_ _0286_ _3428_ _0313_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_5093_ _3528_ _3482_ as2650.r0\[0\] _1206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__4438__A1 _3437_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_797 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4044_ _3561_ _3572_ _3577_ _3443_ _3578_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__7259__CLK clknet_leaf_50_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_83_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5995_ _1909_ _2002_ _2011_ _1104_ _2012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__3749__I _3284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XPHY_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_24_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4946_ _1059_ _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4610__A1 as2650.stack\[3\]\[9\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4877_ _0476_ _0948_ _0993_ _0994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_138_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6616_ as2650.stack\[7\]\[7\] _2603_ _2607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6363__A1 _2130_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3828_ _3240_ _3363_ _3364_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5166__A2 _3372_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6547_ _1288_ _2461_ _2549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3716__A3 _3251_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_118_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_3759_ _3294_ _3295_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XANTENNA__4913__A2 _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_106_503 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6115__A1 _0711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_845 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6478_ _2481_ _2483_ _2484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__5469__A3 _1518_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5429_ _1480_ _1484_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_79_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4677__A1 _0817_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_99_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_43_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_59_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_47_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_25_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_177 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_59_199 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7091__A2 _1066_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_24 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3652__A2 _3184_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1004 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output21_I net21 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5929__A1 as2650.pc\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_394 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3659__I _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_43_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4601__A1 _0718_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5874__I _0664_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_1357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_32_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_10 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5095__B as2650.r0\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_32_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1032 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6106__A1 as2650.stack\[3\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__B2 as2650.stack\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_3_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_140_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6657__A2 _2636_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_729 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_399 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_103 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_412 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_120_583 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3891__A2 _3367_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A1 _3528_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4953__I _0893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_1161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_670 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_372 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_73_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2180 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4800_ _3189_ _0894_ _0922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_61_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5780_ _0663_ _1806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_72_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2191 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6593__A1 _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6593__B2 _2577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4731_ _0827_ _0854_ _0856_ _0077_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_30_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_124_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6345__A1 _2003_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5148__A2 _1246_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4662_ _0807_ _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_119_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6401_ _1885_ _2378_ _1935_ _2409_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_3613_ as2650.cycle\[1\] _3148_ _3149_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_7381_ _0192_ clknet_leaf_30_wb_clk_i as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_134_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4593_ _0702_ _0760_ _0764_ _0031_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_31_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_823 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6332_ _2339_ _2340_ _2341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_115_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_115_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_143_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_131_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6263_ _1963_ _2273_ _2274_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_116_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_837 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__C _1312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5214_ _1324_ _0672_ _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_69_420 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_431 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6194_ as2650.stack\[3\]\[6\] _2206_ _0781_ as2650.stack\[1\]\[6\] _2207_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_135_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_96_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5145_ _1144_ _1257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_637 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7073__A2 _3030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5076_ _0514_ _0578_ _1189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_56_147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6281__B1 _2084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6820__A2 _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4027_ _3528_ _3313_ _3315_ _3560_ _3561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__4831__A1 _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA_clkbuf_leaf_50_wb_clk_i_I clknet_3_5_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6584__A1 _2574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5387__A2 _1133_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5978_ _1439_ _1995_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_100_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4929_ _0675_ _3203_ _1043_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_100_44 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_20_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_60_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_609 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_683 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4103__I _3406_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_182 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7424__CLK clknet_leaf_15_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1287 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_163 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_134_697 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_550 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_699 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3873__A2 _3402_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7064__A2 _3022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A1 as2650.psl\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_29_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_47_158 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_91_916 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_21_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_16_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_62_139 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_44_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_364 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_70_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6575__A1 _1117_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5378__A2 _1284_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_695 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_1080 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_12_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__A1 _2306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6327__B2 _2215_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_11_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6878__A2 _2854_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_89_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4889__A1 _0463_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5550__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_504 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_656 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_537 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_548 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_559 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5853__A3 _1341_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_26_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3864__A2 _3245_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__7055__A2 _2992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_380 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5066__A1 _1060_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_765 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_96_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6802__A2 _2721_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6950_ _2922_ _2923_ _2924_ _2925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or3_1
XFILLER_19_350 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4813__A1 _3451_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5901_ as2650.stack_ptr\[2\] _0648_ _1920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xnor2_1
X_6881_ net32 net51 _2792_ _2859_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_35_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_90_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6015__B1 _1976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_62_662 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_5832_ _1739_ _1675_ _1849_ _1852_ _1853_ _0181_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_50_813 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6566__A1 _1741_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5369__A2 _3151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5763_ _1787_ _1788_ _1789_ _1790_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_37_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4041__A2 _3460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4714_ _0837_ _0845_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_5694_ _0458_ _1725_ _1701_ _1726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_136_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7447__CLK clknet_leaf_53_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7433_ _0244_ clknet_leaf_3_wb_clk_i as2650.r123\[0\]\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_970 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4645_ _0797_ _0050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5019__I _1123_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_119 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7364_ _0175_ clknet_leaf_16_wb_clk_i as2650.cycle\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__4344__A3 _0417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4576_ _0749_ _0736_ _0750_ _0028_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_144_951 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6315_ _2066_ _2318_ _2324_ _1310_ _2325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_116_664 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4858__I _0346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7295_ _0106_ clknet_leaf_44_wb_clk_i as2650.stack\[6\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_143_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_1036 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6246_ _2229_ _2249_ _2257_ _2211_ _2258_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_118_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__B1 _0682_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6177_ _2187_ _2188_ _2189_ _2190_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_57_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_112_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_58_957 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7046__A2 _0419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5128_ _1240_ _1241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A1 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_57_478 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2905 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5059_ _1160_ _1162_ _1164_ _1171_ _1172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_2
XANTENNA__3607__A2 _3142_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2916 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2927 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4804__A1 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_437 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2938 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2949 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4280__A2 _0396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A1 _1764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_71_36 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_55_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_98 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3937__I _3471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4032__A2 _3564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6309__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_138_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_907 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_653 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_973 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_84_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3672__I _3162_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_483 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
Xclkbuf_leaf_36_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_36_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_121_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5296__A1 _0999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_110_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_110_829 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5835__A3 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_423 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_743 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7037__A2 _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5599__A2 _1156_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6796__A1 _2769_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6260__A3 _2098_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_17_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_72_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4271__A2 _0449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_45_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4008__I _3541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_44_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_1175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6548__A1 _3432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_1017 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_38_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4023__A2 _3556_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_211 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_34_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_129_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_61_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_32_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4430_ _0437_ _0597_ _0625_ _0626_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_126_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4326__A3 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4678__I _0717_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4361_ _0557_ _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__inv_1
XFILLER_98_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6100_ _2013_ _2113_ _2114_ _2020_ _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_98_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_623 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_7080_ _1466_ _3035_ _3036_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4292_ _3324_ _0489_ _0490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_98_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_976 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_323 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_133 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6031_ _0699_ _3539_ _2047_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XTAP_345 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5826__A3 _1847_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_356 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_86_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_45_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_367 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5039__A1 _3175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_82_702 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_54_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_724 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_82_757 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6933_ _1891_ _2879_ _2881_ _2909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XPHY_18 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_29 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_278 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6864_ _2173_ _2658_ _2842_ _2843_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_63_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4801__A4 _0875_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_34_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5815_ as2650.cycle\[4\] _1839_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6795_ _1719_ _2633_ _2773_ _2775_ _1763_ _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai221_1
XFILLER_50_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5746_ _1595_ _1773_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_22_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5762__A2 _1490_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__A1 _3308_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5677_ _1711_ _1712_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__5972__I _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7416_ _0227_ clknet_leaf_29_wb_clk_i net35 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_117_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4628_ as2650.stack\[2\]\[1\] _0786_ _0788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6711__A1 net52 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_116_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7347_ _0158_ clknet_leaf_13_wb_clk_i as2650.addr_buff\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_85_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4559_ _0690_ _0737_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_612 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_494 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_334 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7278_ _0089_ clknet_leaf_53_wb_clk_i as2650.psu\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_77_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_678 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_998 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6229_ _2065_ _2240_ _2241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_89_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_54 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3828__A2 _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_65 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_66_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3403 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_862 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3414 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3425 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_100_884 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3436 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3447 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_595 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2702 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3458 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2713 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3469 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_53 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_45_448 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_22_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_234 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_2724 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2735 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2746 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6752__B _3540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4253__A2 _0377_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2757 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_92_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2768 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2779 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3667__I _3202_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_15_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6950__A1 _2922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_127_726 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_51_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_139_597 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_33_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6702__A1 _1807_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5505__A2 _1547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6199__B _2210_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_718 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4498__I _0684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_921 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_965 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5269__A1 _0850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_518 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_0_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_7_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5550__C _1591_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6481__A3 _3382_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_551 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_776 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4492__A2 _3171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6218__I _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_713 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A1 _1242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5122__I _0483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_63_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_532 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5441__A1 _0660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4961__I _1033_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3930_ _3464_ _3465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_45_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3861_ _3395_ _3396_ _3397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_32_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_108_1046 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5600_ _1104_ _1641_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_72_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6580_ _1349_ _2457_ _1583_ _2579_ _2580_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6941__A1 _2151_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3792_ as2650.r123_2\[1\]\[7\] _3328_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6888__I _1683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5531_ _3438_ _1575_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5792__I _1029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_759 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5462_ _1506_ _1514_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7201_ _0012_ clknet_leaf_61_wb_clk_i as2650.r123\[1\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4413_ net8 _0609_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_910 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5393_ _1450_ _1454_ _1455_ _1456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_126_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4201__I _0399_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7132_ _1308_ _3084_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4344_ _0340_ _0321_ _0417_ _0541_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6457__B1 _2460_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7063_ as2650.r123\[0\]\[1\] _3024_ _3026_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4275_ _3300_ _0418_ _0473_ vdd vss gf180mcu_fd_sc_mcu7t5v0__and2_1
XFILLER_80_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_140_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6014_ as2650.stack\[3\]\[2\] _1968_ _1977_ as2650.stack\[2\]\[2\] _2031_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_67_540 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6472__A3 _1168_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A1 _1709_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_132_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_94_370 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_95_893 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5032__I _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_39_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2009 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6224__A3 _2235_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_36_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4235__A2 _0394_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1319 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6916_ _2265_ _2892_ _2893_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6291__C _1886_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6847_ _1348_ _2665_ _2826_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_126_1168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6778_ _2097_ _2758_ _2759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__6932__A1 _1540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_108_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5729_ _1751_ _1756_ _1427_ _1757_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_143_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_136_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5635__C _1576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_578 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_1152 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_64 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_453 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_1049 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_132_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_294 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3200 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_4_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6038__I _2053_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3211 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3222 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_133_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3233 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_381 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3244 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2510 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3255 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_73_554 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3266 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6482__B _0869_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2521 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3277 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2532 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3288 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2543 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3299 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2554 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1820 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2565 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1831 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5974__A2 _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2576 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1842 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2587 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1853 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2598 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3985__A1 _3502_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1864 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1875 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A1 _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_14_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1886 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1897 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__B1 _1298_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_1219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6923__A1 _2000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3737__A1 _3253_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5826__B _1619_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xclkbuf_leaf_51_wb_clk_i clknet_3_5_0_wb_clk_i clknet_leaf_51_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_127_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_108_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6151__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_138_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_123_795 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7100__A1 _3050_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4060_ as2650.holding_reg\[2\] _0261_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_808 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5662__A1 _1637_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_95_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_110_489 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1072 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1045 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_18_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_97_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1078 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A1 _0652_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_51_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_79_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4962_ _1075_ _1076_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__5965__A2 _1938_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_492 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6701_ _3222_ _1811_ _2685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__3976__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3913_ _3296_ _3445_ _3447_ _3448_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
X_4893_ _0569_ _0872_ _1009_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_20_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_33_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6632_ _0665_ _1506_ _1612_ _2617_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
X_3844_ _3318_ _3343_ _3378_ _3379_ _3380_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6914__A1 _2659_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6914__B2 _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3728__A1 _3263_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1010 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6563_ _1218_ _0477_ _2564_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3775_ as2650.r0\[0\] _3311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_118_523 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5193__A3 _0678_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_534 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_34_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5514_ _1557_ _1558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_118_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6494_ _2445_ _2499_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_106_707 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5445_ _1496_ _1497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_133_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_133_526 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_105_217 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_740 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5376_ _0668_ _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__6567__B _2559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7115_ _0466_ _0520_ _3068_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_113_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4327_ _0514_ _0523_ _0524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_101_401 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_141_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7046_ _2993_ _0419_ _3013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_4258_ _0303_ _0455_ _0456_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_102_979 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_27_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4189_ _3246_ _0370_ _0388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_43_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_3_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5697__I _0547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5405__A1 _1466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1105 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_15 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1116 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1127 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5956__A2 _1968_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1149 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7158__A1 _1116_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4106__I _0282_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_10_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_106_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_141_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6905__A1 _2879_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_50_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5708__A2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_810 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6381__A2 _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_52_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_6_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_104_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4392__A1 _3506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_545 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_137_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_342 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_87_1225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_887 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_375 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_74 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6133__A2 _2132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_78_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5892__A1 _0645_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4695__A2 _0828_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_250 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_120_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_78_624 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_732 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_8_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_120_787 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5644__A1 _0862_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_798 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_111_1212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3030 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3041 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3052 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3063 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_73_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3074 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7101__B _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1289 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3085 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_33_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2340 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3096 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2351 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2362 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5947__A2 _1941_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2373 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2384 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1650 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7149__A1 _3319_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2395 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6940__B _2866_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_18_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1661 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1672 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1683 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1694 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7330__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_1196 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_1087 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_31_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3855__I _3390_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_320 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_127_353 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_515 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_142_301 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4135__A1 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5230_ _1082_ _1321_ _1322_ _3434_ _1339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_4
XFILLER_29_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5883__A1 _1488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_529 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_142_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_123_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_38_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_5161_ _3373_ _3548_ _3472_ _3464_ _1273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_123_581 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4112_ _3165_ _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_69_657 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5092_ _1204_ _1205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_64_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5635__A1 _1662_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4438__A2 _0629_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__B1 _2811_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_1129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4043_ _3573_ _3576_ _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_77_690 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_25_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_822 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_40_wb_clk_i_I clknet_3_7_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5994_ _1890_ _2006_ _2008_ _2010_ _2011_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai22_1
XFILLER_36_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4945_ _0677_ _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4610__A2 _0774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4876_ _0500_ _0903_ _0992_ _0929_ _0993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_123_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_18_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6615_ _0721_ _2602_ _2606_ _0211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
X_3827_ _3154_ _3358_ _3362_ _3363_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XANTENNA__7384__D _0195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_128 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_105_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_119_854 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6546_ _0477_ _1854_ _2548_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_119_865 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_10_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3758_ as2650.r0\[0\] _3291_ _3292_ _3293_ as2650.ins_reg\[0\] _3131_ _3294_ vdd
+ vss gf180mcu_fd_sc_mcu7t5v0__mux4_1
XFILLER_134_802 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6477_ _1123_ _2482_ _1520_ _0658_ _2483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XANTENNA__6115__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5980__I _1799_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3689_ _3224_ _3142_ _3225_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_5428_ _1483_ _0147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5469__A4 _1520_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_507 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_0_804 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4596__I _0759_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_710 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_114_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5359_ _1421_ _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_87_410 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_721 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_58_59 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7203__CLK clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5626__A1 _1417_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4429__A2 _0620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_75_616 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7029_ _2988_ _3000_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_21_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_74_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_649 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__6744__C _2726_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3652__A3 _3187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_28_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_15_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_70_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5220__I _1329_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5929__A2 net2 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4264__C _0312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6051__A1 as2650.pc\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_1038 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_output14_I net14 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_19_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_46 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_142_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_11_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_128_117 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_23_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6354__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_7_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_1071 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_137_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_104_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_125_835 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5890__I _1908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6106__A2 _2075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_207 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_827 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_708 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4668__A2 _0810_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5865__A1 _0864_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_719 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_97_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_133_890 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_61_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_592 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_432 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_78_476 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_318 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_627 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5617__A1 _3316_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5093__A2 _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_111_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_59_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_1015 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_1184 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_384 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_46_395 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_61_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2170 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2181 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6670__B _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_37_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2192 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_376 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6593__A2 _1837_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4730_ as2650.stack\[0\]\[9\] _0855_ _0856_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_1480 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1491 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4661_ _0808_ _0809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XANTENNA__6345__A2 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6400_ _1801_ _2407_ _2408_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3612_ as2650.cycle\[0\] _3148_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
X_7380_ _0191_ clknet_leaf_30_wb_clk_i as2650.pc\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4592_ as2650.stack\[3\]\[2\] _0761_ _0764_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_128_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6896__I _1459_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6331_ as2650.pc\[9\] as2650.pc\[8\] _2263_ _2340_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_127_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_183 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA_clkbuf_leaf_7_wb_clk_i_I clknet_3_1_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6262_ _2266_ _2272_ _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_116_879 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7226__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4659__A2 _0806_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_378 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5213_ _0675_ _1324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_175 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_849 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_88_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6193_ _1967_ _2206_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_97_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_443 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5144_ _1183_ _0597_ _1198_ _1076_ _1256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__5608__A1 _0683_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_56_115 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5075_ as2650.psl\[1\] _0579_ _1188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__7376__CLK clknet_leaf_25_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_84_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6564__C _1232_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5084__A2 _1195_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6281__A1 as2650.stack\[1\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4026_ _3450_ _3529_ _3559_ _3484_ _3560_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6281__B2 as2650.stack\[0\]\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_77_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_71_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_65_682 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_991 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_52_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5040__I _1146_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_1542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_94_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4044__B1 _3577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6580__B _1583_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5977_ _1991_ _1993_ _1994_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XANTENNA__5387__A3 _0673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_696 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4595__A1 _0706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_100_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_905 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4928_ _3333_ _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_142_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_90_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_51_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4812__C _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1093 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4859_ _3363_ _0874_ _0977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_138_459 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_5_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_150 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_172 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6529_ _2447_ _0315_ _2516_ _2531_ _2532_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_101_1255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_846 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_69_14 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_107_868 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_49_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A1 _1059_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_326 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5215__I _1325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_667 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_130_860 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_48_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_85_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5862__A4 _1880_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_87_262 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_562 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_882 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_1097 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_435 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_47_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6272__A1 _0729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5075__A2 _0579_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_906 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_608 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_619 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_91_928 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_5_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_939 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_44_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_71_630 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_55_192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6024__A1 _0702_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_71_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_404 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1008 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_138_960 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7249__CLK clknet_leaf_40_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_109_161 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_140_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A1 _1797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_698 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_140_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_516 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_124_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_646 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5125__I _3466_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_337 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_538 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_94_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_117_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_711 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_79_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_1126 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6263__A1 _1963_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5066__A2 _1178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_799 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_90 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4813__A2 _0903_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5900_ _1142_ _1096_ _1919_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_6880_ net33 _2858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_34_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_950 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5831_ _1115_ _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_61_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5369__A3 _0672_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5762_ _1149_ _1490_ _1767_ _1789_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_61_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_6_wb_clk_i clknet_3_1_0_wb_clk_i clknet_leaf_6_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
X_4713_ _0815_ _0838_ _0844_ _0071_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_124_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_5693_ _1235_ _1567_ _1098_ _1725_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6318__A2 _2164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_33_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4329__A1 _3259_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4204__I _0370_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_136_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7432_ _0243_ clknet_leaf_4_wb_clk_i as2650.r123\[0\]\[4\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_15_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4644_ _0731_ as2650.stack\[2\]\[8\] _0784_ _0797_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_141_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7363_ _0174_ clknet_leaf_52_wb_clk_i as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4575_ as2650.stack\[4\]\[12\] _0737_ _0750_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6314_ _2319_ _2320_ _2323_ _1780_ _2324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_7294_ _0105_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_505 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_676 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__5829__A1 _1654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6245_ _2250_ _2251_ _2256_ _1922_ _2257_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_89_549 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__A1 _0666_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6176_ _2187_ _2188_ _2151_ _2189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_69_240 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4501__B2 _0305_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6575__B _2561_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5127_ _1239_ _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_84_210 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_29_137 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_22_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6254__A1 as2650.pc\[8\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5057__A2 _1169_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5058_ _1165_ _1167_ _1170_ _1171_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_84_265 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2906 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2917 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4804__A2 _0925_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2928 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4009_ _3542_ _3543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XTAP_2939 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_129_1100 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_129_1111 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3863__I0 as2650.holding_reg\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4280__A3 _0403_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_25_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6557__A2 _0475_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5765__B1 _1778_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_735 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_90_1276 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XANTENNA__6309__A2 _2312_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3918__I1 as2650.r123_2\[1\]\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6190__B1 _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_621 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3953__I _3442_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_4_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1003 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_1014 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_1074 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_101 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_186 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6493__A1 _3483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_679 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_118_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_49_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_88_571 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_871 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7160__I _3107_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_102_392 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_75_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6245__B2 _1922_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_405 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_416 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6796__A2 _2776_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_112_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_16_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_268 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_91_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6548__A2 _2461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_108_1239 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_125_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_8_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_418 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6720__A2 _3491_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_952 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6379__C _2233_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_126_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4360_ net7 _0557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4731__A1 _0827_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_462 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_98_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_113_613 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_635 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4291_ as2650.r123_2\[0\]\[6\] _0489_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XTAP_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_99_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_98_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6030_ as2650.pc\[2\] net3 _2046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XTAP_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6484__A1 _2468_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_346 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_307 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_input5_I io_in[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_487 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_368 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1070 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_20_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XTAP_379 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_117_1081 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__7070__I _3023_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_221 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_530 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6236__A1 _1307_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5039__A2 _3357_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_541 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_66_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_714 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_574 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6787__A2 _2767_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_224 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6932_ _1540_ _2907_ _2908_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_35_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_19 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_81_257 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7414__CLK clknet_leaf_29_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6863_ _2836_ _2841_ _1689_ _2842_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_62_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5814_ _1797_ _3268_ _1827_ _1838_ _1798_ _0178_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_23_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_6794_ _2633_ _2774_ _2775_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_37_1060 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_52_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5745_ _1740_ _1771_ _1772_ _0175_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_124_1052 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_919 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4970__A1 _1082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3773__A2 _3241_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_124_1085 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5676_ _1241_ _1266_ _1711_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_727 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_135_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7415_ _0226_ clknet_leaf_29_wb_clk_i net34 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XANTENNA__7392__D _0203_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4627_ _0647_ _0785_ _0787_ _0042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XANTENNA__6711__A2 _2654_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_117_963 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_11_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4558_ _0691_ _0736_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7346_ _0157_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_104_602 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_117_996 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_144_782 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_324 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_944 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_81_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_7277_ _0088_ clknet_leaf_6_wb_clk_i as2650.r123_2\[2\]\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4489_ _3197_ _0676_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_2
XFILLER_106_11 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_22 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6475__A1 _1506_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_988 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6228_ _2230_ _2232_ _2239_ _1310_ _2240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
XFILLER_77_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_103_178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_58_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_26 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6159_ _0718_ _1984_ _2172_ _0189_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_131_1023 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_891 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3404 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3415 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_874 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3426 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3437 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3448 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2703 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2714 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3459 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4789__A1 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2725 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2736 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2747 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5450__A2 _1501_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4253__A3 _0450_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2758 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2769 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5649__B _1687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_53_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_53_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3948__I _3482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_13_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5202__A2 _1264_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1040 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_90_1051 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_40_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_543 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A2 _2923_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_107_1261 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1272 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_16_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_127_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_1283 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_1147 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_31_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6702__A2 _2660_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_120_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_68_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6199__C _2211_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_107_473 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_270 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_68_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput40 net40 io_out[3] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XANTENNA__6466__A1 _1132_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_110_605 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_95_338 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_95_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5403__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_48_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7437__CLK clknet_leaf_52_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_1216 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_76_585 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6769__A2 _2191_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4019__I _3552_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_17_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_63_246 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_44_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3860_ _3161_ _3208_ _3396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__4182__C _0300_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_72_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_3791_ _3326_ _3327_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_108_1069 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6941__A2 _2906_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_34_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XPHY_190 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_121_1203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_9_851 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5530_ net21 _1571_ _1574_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_117_215 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5461_ _1512_ _1513_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_51_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7200_ _0011_ clknet_leaf_63_wb_clk_i as2650.r123\[1\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4412_ _3366_ _0607_ _0608_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
X_5392_ _3204_ _1455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_114_900 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_933 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7131_ _1572_ _0579_ _3083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4343_ _0538_ _0539_ _0540_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_2
XFILLER_98_110 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_67_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_98_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_421 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_655 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_99_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_966 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_59_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7062_ _3437_ _3022_ _3025_ _0239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_99_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_115_1007 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4274_ _0320_ _0471_ _0472_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_115_1018 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_98_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_45_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_80_1231 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6013_ _1920_ _2030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_101_638 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7014__B _1620_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6409__I _2415_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6472__A4 _1657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6209__A1 _0720_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5680__A2 _1713_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1309 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_82_566 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5432__A2 _1477_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_717 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6915_ _2267_ _2817_ _2269_ _2892_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_82_599 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_63_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_74_1024 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_62_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6846_ _1272_ _0568_ _2824_ _2825_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor3_1
XFILLER_126_1136 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_50_452 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5196__A1 _1042_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6393__B1 _0754_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6777_ _2043_ _2757_ _2758_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__5983__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_22_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_3989_ _3523_ _3524_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_17_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4943__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5916__C _1853_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5728_ _1649_ _1754_ _1755_ _1756_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_108_226 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5659_ _1695_ _3434_ _1696_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_108_237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_85_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_730 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_43 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7329_ _0140_ clknet_leaf_25_wb_clk_i as2650.stack_ptr\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_116_292 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_121 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_903 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_977 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_132_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_76 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_914 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_77_47 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_105_999 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_28_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_131_273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_498 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5120__A1 _1231_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5223__I _1238_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_58_552 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5671__A2 _1706_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_3201 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3212 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA_output44_I net44 vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_85_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_100_671 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3223 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3234 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_46_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_3245 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_85_393 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2500 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3256 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_22_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2511 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3267 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2522 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2533 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3278 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3289 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2544 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_60_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1810 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2555 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3678__I _3213_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1821 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_92_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_2566 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1832 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2577 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1843 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2588 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1854 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_53_290 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_42_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__3985__A2 _3355_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2599 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_1865 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1876 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__7176__A2 _1729_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1887 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1898 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__5187__A1 as2650.psu\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5187__B2 as2650.psu\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_35_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__3737__A2 _3256_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_373 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4302__I _0342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_218 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5842__B _3237_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_1237 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_925 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_1_570 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_68_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_122_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_66 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_7_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_77_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5662__A2 _1698_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_91 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_3_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_76_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA_clkbuf_leaf_30_wb_clk_i_I clknet_3_6_0_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_64_544 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1057 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_92_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6611__A1 _0710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_352 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5414__A2 _1457_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_92_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4961_ _1033_ _1075_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_45_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_396 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6700_ _2648_ _2684_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_75_1344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3912_ _3367_ _3446_ _3388_ _3447_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
X_4892_ _0546_ _0878_ _0945_ _1007_ _1008_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_32_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_6631_ _1558_ _2615_ _2616_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3843_ _3312_ _3379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__3728__A2 _3242_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4925__A1 _1034_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_20_669 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_3774_ _3309_ _3310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_6562_ _1296_ _1092_ _2562_ _2563_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_121_1022 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6390__A3 _2397_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5193__A4 _1108_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_121_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7009__B _1461_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5513_ _0661_ _3359_ _1557_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_6493_ _3483_ _2497_ _2498_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_118_557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_118_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5444_ _3215_ _3216_ _3218_ as2650.cycle\[0\] _1496_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_2
XFILLER_12_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_105_229 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4153__A2 _0332_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5350__A1 _0858_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5375_ _1429_ _1431_ _1432_ _1437_ _1438_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XFILLER_82_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6567__C _2567_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_114_763 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7114_ _0445_ _0974_ _0466_ _0520_ _3067_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi22_1
X_4326_ _0374_ _0377_ _0450_ _0522_ _0523_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XFILLER_101_413 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_796 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5102__A1 _1173_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7045_ net42 _3012_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XFILLER_59_349 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4257_ _3259_ _0449_ _0454_ _0455_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_102_969 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_113_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_446 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6850__A1 _1100_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_86_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4188_ as2650.holding_reg\[4\] _0262_ _0387_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_132_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5978__I _1439_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_67_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6583__B _2569_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_28_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_330 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_23_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_56 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_82_363 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5199__B _1310_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6602__A1 as2650.stack\[7\]\[1\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_728 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_1106 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1117 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_63_27 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_103_78 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1128 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_93_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1139 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_70_547 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_70_558 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5927__B _1422_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5169__A1 as2650.psl\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6829_ _1689_ _2808_ _2809_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_51_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4831__B _0917_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_23_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_143_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_844 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_136_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_10_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_136_332 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_104_1286 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_30_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_109_579 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_13 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7282__CLK clknet_leaf_60_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5662__B _1097_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_97 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3961__I _3435_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_105_752 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_68 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_700 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5892__A2 _1889_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_65_1557 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_2_389 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_52 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6049__I _1525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_104_295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_606 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_120_777 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_77_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_617 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_4_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_92_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_980 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_691 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3020 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3031 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3042 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3053 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_74_875 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_98_1377 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3064 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3075 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2330 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3086 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2341 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_27_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2352 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_3097 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2363 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2374 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1640 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3958__A2 _3492_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2385 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1651 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__4080__A1 as2650.holding_reg\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2396 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_109_1120 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_1662 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1673 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_72_1528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_144_1033 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_14_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_109_1153 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_1684 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1695 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__6357__B1 _0805_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_144_1077 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6512__I _1201_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_70_1241 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_811 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5580__A1 _3209_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_866 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5128__I _1240_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_128_899 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_115_527 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_6_673 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_127_398 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4967__I as2650.halted vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_143_869 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_68_1170 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5883__A2 _3293_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5160_ _1212_ _1272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_116_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_69_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_116_1113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__3894__A1 _3398_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4111_ _0292_ _0301_ _0304_ _0309_ _0310_ _0311_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai32_2
XANTENNA__7085__A1 _1046_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_97_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5091_ _1203_ _1204_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_110_232 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_68_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_96_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_110_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_111_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5635__A2 _1673_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6832__A1 _2141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4042_ _3574_ _3568_ _3575_ _3576_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_2
XANTENNA__6832__B2 _1428_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_68_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3646__A1 _3180_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_49_371 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_83_127 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_110_298 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_83_149 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_374 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5399__A1 _0751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_91_160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5993_ _2009_ _1994_ _2010_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XANTENNA__4207__I _0405_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4944_ _1041_ _1057_ _1058_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4071__A1 _3419_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_80_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_33_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4875_ _0989_ _0915_ _0962_ _0991_ _0992_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
XFILLER_60_591 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6614_ as2650.stack\[7\]\[6\] _2603_ _2606_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3826_ _3361_ _3362_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_21_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_119_833 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_321 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5571__A1 _3214_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6545_ _0422_ _1837_ _2547_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_3757_ as2650.r123\[2\]\[0\] as2650.r123_2\[2\]\[0\] as2650.psl\[4\] _3293_ vdd vss
+ gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_134_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_302 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_6476_ _1502_ _2482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_3688_ as2650.cycle\[7\] _3224_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_9 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5427_ as2650.r123_2\[0\]\[4\] _0987_ _1480_ _1483_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XANTENNA__4126__A2 _0325_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5323__A1 as2650.stack\[5\]\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_133_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_519 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_260 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5358_ _1336_ _0671_ _1421_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_114_582 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_1156 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_956 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_733 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7076__A1 _0572_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_59_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4309_ _3309_ _0502_ _0506_ _0507_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_82_1178 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_744 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_455 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5289_ as2650.r123_2\[1\]\[2\] _0958_ _1378_ _1379_ vdd vss gf180mcu_fd_sc_mcu7t5v0__mux2_2
XFILLER_101_243 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_102_766 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5626__A2 _0657_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6823__A1 _0482_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_74_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_7028_ _3483_ _2996_ _2998_ _2999_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi21_1
XFILLER_60_1454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_74_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5501__I _1535_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_56_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_83_672 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_70_300 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6051__A2 _2001_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_128_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4117__I _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_70_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_58_1383 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_87 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_93_1274 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_24_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1304 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_93_1296 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_141_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_15_1209 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_135_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_71_1561 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_128_129 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4365__A2 _0550_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5562__A1 _1069_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_137_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_11_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_104_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_85 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_663 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_109_354 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_125_814 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_136_151 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_1034 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_109_387 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_125_847 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_139_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_87_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_89 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_195 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_69_1490 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_97_219 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5865__A2 _1613_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_140_839 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_117_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__3876__A1 as2650.psl\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_79_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_94_915 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_926 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5617__A2 _1155_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6814__A1 _1269_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_78_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_66_639 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3628__A1 _3161_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_93_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5093__A3 as2650.r0\[0\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_111_1021 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_24_1095 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_0_1009 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_80_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6951__B _2715_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_61_311 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6578__B1 _0549_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_94_1027 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6042__A2 _2014_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2160 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_76_1450 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2171 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_61_366 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_62_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2182 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_21_208 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2193 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_1470 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_15_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_1481 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XANTENNA__3800__A1 _3194_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_1492 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_119_107 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4660_ _0807_ _0808_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_3611_ _3146_ _3147_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_4591_ _0697_ _0760_ _0763_ _0030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_116_803 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
X_6330_ as2650.pc\[10\] _2339_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_7_993 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_50_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_644 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__4108__A2 _0306_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_115_335 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6261_ _2269_ _2271_ _2272_ vdd vss gf180mcu_fd_sc_mcu7t5v0__or2_1
XFILLER_89_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_115_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_103_508 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5212_ _0610_ _1126_ _1323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XANTENNA__7006__C _2432_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_69_400 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_130_327 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_880 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_97_720 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6192_ _2203_ _2204_ _2205_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_142_187 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5143_ _1254_ _1255_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkinv_1
XANTENNA__6618__S _2595_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_9_1067 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5608__A2 _0685_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_131_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_403 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_56_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5074_ _0394_ _0467_ _0536_ _1186_ _1187_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor4_1
XFILLER_69_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_96_285 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_56_138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_42_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4025_ _3452_ _3537_ _3558_ _3479_ _3559_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai211_1
XANTENNA__6281__A2 _2082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5321__I _1396_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__4292__A1 _3324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_38_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_65_661 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_65_694 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_80_620 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_92_480 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_80_642 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_129_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_52_355 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_13_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5976_ _1946_ _1947_ _1992_ _1993_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_80_686 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5387__A4 _1449_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4927_ _1030_ _1040_ _1041_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__4595__A2 _0760_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_127_1061 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_4858_ _0346_ _0976_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_53_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5544__A1 _1577_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_3809_ _3344_ _3345_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__4347__A2 _0543_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_119_641 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
X_4789_ _3302_ _0873_ _0909_ _0910_ _0911_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi211_1
X_6528_ _2499_ _2529_ _2530_ _2531_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_107_825 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_313 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1267 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_6 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6101__B _2115_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6459_ _1088_ _2465_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_109_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_134_666 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_357 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_109_99 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_136_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_828 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5847__A2 _1064_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__3858__A1 _3302_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_88_742 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_87_230 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__7320__CLK clknet_leaf_42_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_134_1054 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_75_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_21_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_69 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_28_385 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6024__A2 _1984_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_344 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_44_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_70_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4035__A1 _3388_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_71_675 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_19_1131 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5783__A1 _1639_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_54_1099 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_7_212 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_89_1118 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_994 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_137_471 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_611 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_32_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_137_482 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_124_132 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_124_143 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XFILLER_113_817 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5838__A2 _3141_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_98_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_506 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_517 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_26_1102 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_528 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_79_731 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XTAP_539 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_59_70 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_850 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_121_861 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_78_263 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_360 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_94_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_734 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_120_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_436 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_113_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_66_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6263__A2 _2273_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_43_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_93_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_93_266 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4274__A1 _0320_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_81_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_75_80 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_940 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6015__A2 _2025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5830_ _1739_ _1620_ _1851_ _1852_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor3_1
XFILLER_61_130 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_50_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5761_ _1778_ _1762_ _1768_ _1788_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__3596__I _3131_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4712_ as2650.stack\[0\]\[3\] _0839_ _0844_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_72_1166 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5692_ _1724_ _0170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
X_7431_ _0242_ clknet_leaf_63_wb_clk_i as2650.r123\[0\]\[3\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_120_1109 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4329__A2 _0525_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_4643_ _0726_ _0791_ _0796_ _0049_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_102_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_11_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6700__I _2648_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_983 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_128_460 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7362_ _0173_ clknet_leaf_7_wb_clk_i as2650.holding_reg\[7\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
X_4574_ _0748_ _0749_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_116_633 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_102_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6313_ _1959_ _2322_ _2323_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_144_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_7293_ _0104_ clknet_leaf_43_wb_clk_i as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_131_603 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4220__I _0418_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5829__A2 _1850_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_118_1016 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_103_305 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6244_ as2650.stack\[1\]\[7\] _2252_ _2253_ as2650.stack\[0\]\[7\] _2255_ _2256_
+ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_103_316 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_143_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6856__B _2834_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_124 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_115_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_130_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__4501__A2 _0667_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_6175_ _0558_ _0486_ _2188_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_130_157 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4501__B3 _0687_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_130_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_85_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_130_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_112_883 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_5126_ _3538_ _1239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_84_200 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_111_382 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6254__A2 _0558_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_84_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_84_244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_73_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5057_ _1168_ _1169_ _3152_ _1170_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XTAP_2907 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_44_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2918 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_4008_ _3541_ _3542_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XTAP_2929 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5986__I as2650.addr_buff\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__6006__A2 _2022_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_1134 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_38_1028 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_26_889 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__4017__A1 _3346_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_40_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_111_67 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5765__A1 _1030_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1222 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_5959_ _0753_ _1977_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XANTENNA__5765__B2 _1781_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_1233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_142_1312 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_139_703 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_16_1315 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_90_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_51_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_138_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_747 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5517__A1 _0920_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5427__S _1480_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_5_705 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_101_1020 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__5654__C _1691_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_931 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6190__B2 as2650.stack\[6\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_101_1042 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_88_1173 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_101_1064 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_49_1135 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_134_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_154 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_107_677 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_688 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_1_922 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_106_176 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_121_113 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__6766__B _2747_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_122_647 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_106_198 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_27_1422 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__6493__A2 _2497_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_0_454 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_88_594 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_62_1379 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_29_73 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_48_447 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_48_469 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_75_255 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_76_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_5_1273 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_112_1160 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_63_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_99_1280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_225 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_95_1122 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_99_1291 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5896__I _1914_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_90_247 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_43_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_32_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xclkbuf_leaf_45_wb_clk_i clknet_3_7_0_wb_clk_i clknet_leaf_45_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XFILLER_71_472 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7216__CLK clknet_leaf_33_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XANTENNA__5756__A1 _1779_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_73_1486 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_84_8 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_909 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__7366__CLK clknet_leaf_14_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_129_279 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6181__A1 _2007_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_8_598 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_144_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_1202 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_126_975 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_99_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5136__I _3152_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_125_485 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4290_ as2650.r0\[6\] _3199_ _0488_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XTAP_303 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_84_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_113_658 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_140_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_325 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_146 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_347 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_358 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_112_168 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_67_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_369 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_67_723 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_112_179 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_132_1525 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_121_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_41_1419 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_39_425 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__6236__A2 _2013_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_13_2 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__5039__A3 _1150_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_55_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_67_778 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_26_108 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_66_277 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_94_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6931_ _1891_ _2885_ _2887_ _2907_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_54_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5995__A1 _1909_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_66_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_81_236 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6862_ _2173_ _2837_ _2840_ _2644_ _1257_ _2841_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_81_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_78_1386 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_39_1348 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_90_770 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5813_ _1830_ _1835_ _1836_ _1837_ _1577_ _1838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__aoi221_1
XFILLER_22_314 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6793_ _2770_ _2772_ _2771_ _2774_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_91_1564 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_5744_ _1575_ _1772_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
XFILLER_124_1031 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__4970__A2 _1083_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5675_ _3528_ _1710_ vdd vss gf180mcu_fd_sc_mcu7t5v0__buf_1
X_7414_ _0225_ clknet_leaf_29_wb_clk_i net33 vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_129_780 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4626_ as2650.stack\[2\]\[0\] _0786_ _0787_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XFILLER_102_1340 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_430 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7345_ _0156_ clknet_leaf_12_wb_clk_i as2650.addr_buff\[5\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_89_1493 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_4557_ _0734_ _0735_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_144_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_116_463 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_614 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_46_1308 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_104_625 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_7276_ _0087_ clknet_leaf_62_wb_clk_i as2650.r123_2\[2\]\[6\] vdd vss gf180mcu_fd_sc_mcu7t5v0__dffq_1
XFILLER_143_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_89_336 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4488_ _3206_ _0675_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_131_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_6227_ _2236_ _2238_ _2239_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
XANTENNA__6475__A2 _1342_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_106_34 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_131_488 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_131_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_98_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_870 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_6158_ _2130_ _2171_ _2039_ _2172_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_112_680 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_131_1013 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_881 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_892 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_100_842 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_85_542 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_3405 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
X_5109_ _1220_ _3342_ _0553_ _1221_ _1222_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai31_1
XTAP_3416 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_6_1560 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
X_6089_ _0704_ _2067_ _2104_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_2
XFILLER_58_789 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XTAP_3427 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_417 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_886 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_3438 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_131_1079 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_72_203 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_85_586 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XTAP_3449 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_428 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XANTENNA__7239__CLK clknet_leaf_39_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XTAP_2704 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_45_439 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_57_299 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XTAP_2715 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XTAP_2726 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_2_1457 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XTAP_2737 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_57_1415 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2748 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_122_88 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_60_409 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_72_269 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_82_37 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XTAP_2759 vdd vss gf180mcu_fd_sc_mcu7t5v0__filltie
XFILLER_25_141 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_14_815 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_144_1407 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_92_1339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__5738__A1 _1527_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_41_634 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1181 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_0_1192 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_80_280 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4125__I _0324_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_511 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6950__A3 _2924_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_139_555 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_107_1295 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_139_577 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
Xclkbuf_opt_2_1_wb_clk_i clknet_opt_2_0_wb_clk_i clknet_opt_2_1_wb_clk_i vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_16
XANTENNA__6340__I _2321_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_103_1159 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_126_238 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_108_953 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__4713__A2 _0838_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_135_761 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_135_772 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_135_783 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
Xoutput30 net30 io_out[1] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_135_794 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
Xoutput41 net41 io_out[4] vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_3
XFILLER_107_496 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_122_433 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_122_444 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_123_978 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6466__A2 _3314_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_96_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_32
XFILLER_123_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_49_712 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XANTENNA__7104__C _1785_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_76_531 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_48_233 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_114_1244 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_23_1138 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_37_918 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_97_1206 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_76_575 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_97_1228 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_64_737 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_131_1580 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_63_258 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_91_567 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_72_792 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XANTENNA__5729__A1 _1751_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_31_144 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_20_818 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
X_3790_ _3133_ _3198_ _3326_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nor2_1
XFILLER_125_1351 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_64
XFILLER_82_5 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XPHY_180 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XPHY_191 vdd vss gf180mcu_fd_sc_mcu7t5v0__endcap
XFILLER_117_205 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_118_739 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_12_1521 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
X_5460_ _1493_ _1512_ vdd vss gf180mcu_fd_sc_mcu7t5v0__clkbuf_1
XFILLER_117_227 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_117_249 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_133_709 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_4411_ _3338_ _0606_ _0607_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_2
XFILLER_12_1576 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XANTENNA__5901__A1 as2650.stack_ptr\[2\] vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_5391_ _0658_ _1453_ _0673_ _1454_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_114_912 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_7130_ _1184_ _3071_ _3082_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_114_923 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
X_4342_ _0468_ _0418_ _0525_ _0539_ vdd vss gf180mcu_fd_sc_mcu7t5v0__oai21_1
XFILLER_114_945 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_125_282 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_119_1155 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XANTENNA__6457__A2 _3343_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
X_7061_ as2650.r123\[0\]\[0\] _3024_ _3025_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand2_1
X_4273_ _0470_ _0417_ _0471_ vdd vss gf180mcu_fd_sc_mcu7t5v0__xor2_1
XFILLER_99_689 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_113_466 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_4
XFILLER_114_989 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_306 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_86_317 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_101_628 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_8
XFILLER_86_328 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
X_6012_ _2024_ _2026_ _2028_ _2029_ vdd vss gf180mcu_fd_sc_mcu7t5v0__nand3_1
XFILLER_98_188 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
XFILLER_100_105 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_1
XFILLER_86_339 vdd vss gf180mcu_fd_sc_mcu7t5v0__fillcap_16
XANTENNA__7014__C _1164_ vdd vss gf180mcu_fd_sc_mcu7t5v0__antenna
XFILLER_113_499 vdd vss gf180mcu_fd_sc_mcu7t5v0__fill_2
.ends

