magic
tech gf180mcuD
magscale 1 10
timestamp 1701964274
<< metal1 >>
rect 50418 51886 50430 51938
rect 50482 51935 50494 51938
rect 51650 51935 51662 51938
rect 50482 51889 51662 51935
rect 50482 51886 50494 51889
rect 51650 51886 51662 51889
rect 51714 51886 51726 51938
rect 1344 51770 53648 51804
rect 1344 51718 19838 51770
rect 19890 51718 19942 51770
rect 19994 51718 20046 51770
rect 20098 51718 50558 51770
rect 50610 51718 50662 51770
rect 50714 51718 50766 51770
rect 50818 51718 53648 51770
rect 1344 51684 53648 51718
rect 41246 51602 41298 51614
rect 41246 51538 41298 51550
rect 41470 51602 41522 51614
rect 41470 51538 41522 51550
rect 50542 51602 50594 51614
rect 50542 51538 50594 51550
rect 41794 51438 41806 51490
rect 41858 51438 41870 51490
rect 49982 51378 50034 51390
rect 49982 51314 50034 51326
rect 50430 51378 50482 51390
rect 50430 51314 50482 51326
rect 50654 51378 50706 51390
rect 50654 51314 50706 51326
rect 51214 51378 51266 51390
rect 51214 51314 51266 51326
rect 51438 51378 51490 51390
rect 51438 51314 51490 51326
rect 51662 51378 51714 51390
rect 51662 51314 51714 51326
rect 49758 51266 49810 51278
rect 49758 51202 49810 51214
rect 51326 51266 51378 51278
rect 51326 51202 51378 51214
rect 1344 50986 53648 51020
rect 1344 50934 4478 50986
rect 4530 50934 4582 50986
rect 4634 50934 4686 50986
rect 4738 50934 35198 50986
rect 35250 50934 35302 50986
rect 35354 50934 35406 50986
rect 35458 50934 53648 50986
rect 1344 50900 53648 50934
rect 51102 50818 51154 50830
rect 51102 50754 51154 50766
rect 18498 50654 18510 50706
rect 18562 50654 18574 50706
rect 31042 50654 31054 50706
rect 31106 50654 31118 50706
rect 40338 50654 40350 50706
rect 40402 50654 40414 50706
rect 41234 50654 41246 50706
rect 41298 50654 41310 50706
rect 48290 50654 48302 50706
rect 48354 50654 48366 50706
rect 24334 50594 24386 50606
rect 15698 50542 15710 50594
rect 15762 50542 15774 50594
rect 24334 50530 24386 50542
rect 24782 50594 24834 50606
rect 24782 50530 24834 50542
rect 27134 50594 27186 50606
rect 27134 50530 27186 50542
rect 27694 50594 27746 50606
rect 33954 50542 33966 50594
rect 34018 50542 34030 50594
rect 37426 50542 37438 50594
rect 37490 50542 37502 50594
rect 44146 50542 44158 50594
rect 44210 50542 44222 50594
rect 45490 50542 45502 50594
rect 45554 50542 45566 50594
rect 51650 50542 51662 50594
rect 51714 50542 51726 50594
rect 27694 50530 27746 50542
rect 23998 50482 24050 50494
rect 16370 50430 16382 50482
rect 16434 50430 16446 50482
rect 23998 50418 24050 50430
rect 24110 50482 24162 50494
rect 24110 50418 24162 50430
rect 24558 50482 24610 50494
rect 24558 50418 24610 50430
rect 25006 50482 25058 50494
rect 25006 50418 25058 50430
rect 25118 50482 25170 50494
rect 25118 50418 25170 50430
rect 27358 50482 27410 50494
rect 27358 50418 27410 50430
rect 27582 50482 27634 50494
rect 44942 50482 44994 50494
rect 33170 50430 33182 50482
rect 33234 50430 33246 50482
rect 38210 50430 38222 50482
rect 38274 50430 38286 50482
rect 43362 50430 43374 50482
rect 43426 50430 43438 50482
rect 46162 50430 46174 50482
rect 46226 50430 46238 50482
rect 27582 50418 27634 50430
rect 44942 50418 44994 50430
rect 18958 50370 19010 50382
rect 18958 50306 19010 50318
rect 34414 50370 34466 50382
rect 34414 50306 34466 50318
rect 37102 50370 37154 50382
rect 37102 50306 37154 50318
rect 48750 50370 48802 50382
rect 48750 50306 48802 50318
rect 1344 50202 53648 50236
rect 1344 50150 19838 50202
rect 19890 50150 19942 50202
rect 19994 50150 20046 50202
rect 20098 50150 50558 50202
rect 50610 50150 50662 50202
rect 50714 50150 50766 50202
rect 50818 50150 53648 50202
rect 1344 50116 53648 50150
rect 17726 50034 17778 50046
rect 17726 49970 17778 49982
rect 24110 50034 24162 50046
rect 24110 49970 24162 49982
rect 27582 50034 27634 50046
rect 27582 49970 27634 49982
rect 37774 50034 37826 50046
rect 37774 49970 37826 49982
rect 38446 50034 38498 50046
rect 38446 49970 38498 49982
rect 49646 50034 49698 50046
rect 49646 49970 49698 49982
rect 26910 49922 26962 49934
rect 18498 49870 18510 49922
rect 18562 49870 18574 49922
rect 20738 49870 20750 49922
rect 20802 49870 20814 49922
rect 26910 49858 26962 49870
rect 27358 49922 27410 49934
rect 31054 49922 31106 49934
rect 28578 49870 28590 49922
rect 28642 49870 28654 49922
rect 27358 49858 27410 49870
rect 31054 49858 31106 49870
rect 31950 49922 32002 49934
rect 31950 49858 32002 49870
rect 42030 49922 42082 49934
rect 51090 49870 51102 49922
rect 51154 49870 51166 49922
rect 42030 49858 42082 49870
rect 17390 49810 17442 49822
rect 17390 49746 17442 49758
rect 17726 49810 17778 49822
rect 17726 49746 17778 49758
rect 18062 49810 18114 49822
rect 25454 49810 25506 49822
rect 18722 49758 18734 49810
rect 18786 49758 18798 49810
rect 20066 49758 20078 49810
rect 20130 49758 20142 49810
rect 25218 49758 25230 49810
rect 25282 49758 25294 49810
rect 18062 49746 18114 49758
rect 25454 49746 25506 49758
rect 25678 49810 25730 49822
rect 25678 49746 25730 49758
rect 25790 49810 25842 49822
rect 27246 49810 27298 49822
rect 37438 49810 37490 49822
rect 26450 49758 26462 49810
rect 26514 49758 26526 49810
rect 26674 49758 26686 49810
rect 26738 49758 26750 49810
rect 27906 49758 27918 49810
rect 27970 49758 27982 49810
rect 31266 49758 31278 49810
rect 31330 49758 31342 49810
rect 33954 49758 33966 49810
rect 34018 49758 34030 49810
rect 25790 49746 25842 49758
rect 27246 49746 27298 49758
rect 37438 49746 37490 49758
rect 37550 49810 37602 49822
rect 37550 49746 37602 49758
rect 37886 49810 37938 49822
rect 48750 49810 48802 49822
rect 38658 49758 38670 49810
rect 38722 49758 38734 49810
rect 50306 49758 50318 49810
rect 50370 49758 50382 49810
rect 37886 49746 37938 49758
rect 48750 49746 48802 49758
rect 19630 49698 19682 49710
rect 23214 49698 23266 49710
rect 22866 49646 22878 49698
rect 22930 49646 22942 49698
rect 19630 49634 19682 49646
rect 23214 49634 23266 49646
rect 25566 49698 25618 49710
rect 31726 49698 31778 49710
rect 37662 49698 37714 49710
rect 48302 49698 48354 49710
rect 26786 49646 26798 49698
rect 26850 49646 26862 49698
rect 30706 49646 30718 49698
rect 30770 49646 30782 49698
rect 32050 49646 32062 49698
rect 32114 49646 32126 49698
rect 34738 49646 34750 49698
rect 34802 49646 34814 49698
rect 36866 49646 36878 49698
rect 36930 49646 36942 49698
rect 42130 49646 42142 49698
rect 42194 49646 42206 49698
rect 25566 49634 25618 49646
rect 31726 49634 31778 49646
rect 37662 49634 37714 49646
rect 48302 49634 48354 49646
rect 49198 49698 49250 49710
rect 49198 49634 49250 49646
rect 49982 49698 50034 49710
rect 53218 49646 53230 49698
rect 53282 49646 53294 49698
rect 49982 49634 50034 49646
rect 23438 49586 23490 49598
rect 23438 49522 23490 49534
rect 23662 49586 23714 49598
rect 23662 49522 23714 49534
rect 38334 49586 38386 49598
rect 38334 49522 38386 49534
rect 41806 49586 41858 49598
rect 41806 49522 41858 49534
rect 48974 49586 49026 49598
rect 48974 49522 49026 49534
rect 1344 49418 53648 49452
rect 1344 49366 4478 49418
rect 4530 49366 4582 49418
rect 4634 49366 4686 49418
rect 4738 49366 35198 49418
rect 35250 49366 35302 49418
rect 35354 49366 35406 49418
rect 35458 49366 53648 49418
rect 1344 49332 53648 49366
rect 19294 49250 19346 49262
rect 19294 49186 19346 49198
rect 27134 49250 27186 49262
rect 27134 49186 27186 49198
rect 35086 49250 35138 49262
rect 35086 49186 35138 49198
rect 35422 49250 35474 49262
rect 35422 49186 35474 49198
rect 27246 49138 27298 49150
rect 16370 49086 16382 49138
rect 16434 49086 16446 49138
rect 27246 49074 27298 49086
rect 38334 49138 38386 49150
rect 38334 49074 38386 49086
rect 41246 49138 41298 49150
rect 51886 49138 51938 49150
rect 47058 49086 47070 49138
rect 47122 49086 47134 49138
rect 41246 49074 41298 49086
rect 51886 49074 51938 49086
rect 18174 49026 18226 49038
rect 19966 49026 20018 49038
rect 13570 48974 13582 49026
rect 13634 48974 13646 49026
rect 19618 48974 19630 49026
rect 19682 48974 19694 49026
rect 18174 48962 18226 48974
rect 19966 48962 20018 48974
rect 38222 49026 38274 49038
rect 38222 48962 38274 48974
rect 38558 49026 38610 49038
rect 41134 49026 41186 49038
rect 40898 48974 40910 49026
rect 40962 48974 40974 49026
rect 38558 48962 38610 48974
rect 41134 48962 41186 48974
rect 48750 49026 48802 49038
rect 48750 48962 48802 48974
rect 48974 49026 49026 49038
rect 48974 48962 49026 48974
rect 49198 49026 49250 49038
rect 49746 48974 49758 49026
rect 49810 48974 49822 49026
rect 49198 48962 49250 48974
rect 18398 48914 18450 48926
rect 14242 48862 14254 48914
rect 14306 48862 14318 48914
rect 18398 48850 18450 48862
rect 18510 48914 18562 48926
rect 18510 48850 18562 48862
rect 20302 48914 20354 48926
rect 20302 48850 20354 48862
rect 35198 48914 35250 48926
rect 35198 48850 35250 48862
rect 37998 48914 38050 48926
rect 37998 48850 38050 48862
rect 41358 48914 41410 48926
rect 41358 48850 41410 48862
rect 41582 48914 41634 48926
rect 41582 48850 41634 48862
rect 46734 48914 46786 48926
rect 46734 48850 46786 48862
rect 47182 48914 47234 48926
rect 47182 48850 47234 48862
rect 16830 48802 16882 48814
rect 16830 48738 16882 48750
rect 19406 48802 19458 48814
rect 19406 48738 19458 48750
rect 20190 48802 20242 48814
rect 20190 48738 20242 48750
rect 30942 48802 30994 48814
rect 30942 48738 30994 48750
rect 37102 48802 37154 48814
rect 37102 48738 37154 48750
rect 38446 48802 38498 48814
rect 38446 48738 38498 48750
rect 46398 48802 46450 48814
rect 46398 48738 46450 48750
rect 46958 48802 47010 48814
rect 46958 48738 47010 48750
rect 48302 48802 48354 48814
rect 48302 48738 48354 48750
rect 1344 48634 53648 48668
rect 1344 48582 19838 48634
rect 19890 48582 19942 48634
rect 19994 48582 20046 48634
rect 20098 48582 50558 48634
rect 50610 48582 50662 48634
rect 50714 48582 50766 48634
rect 50818 48582 53648 48634
rect 1344 48548 53648 48582
rect 21534 48466 21586 48478
rect 21534 48402 21586 48414
rect 22206 48466 22258 48478
rect 22206 48402 22258 48414
rect 25678 48466 25730 48478
rect 25678 48402 25730 48414
rect 27022 48466 27074 48478
rect 27022 48402 27074 48414
rect 27134 48466 27186 48478
rect 46846 48466 46898 48478
rect 39778 48414 39790 48466
rect 39842 48414 39854 48466
rect 42130 48414 42142 48466
rect 42194 48414 42206 48466
rect 27134 48402 27186 48414
rect 46846 48402 46898 48414
rect 49982 48466 50034 48478
rect 49982 48402 50034 48414
rect 50206 48466 50258 48478
rect 50206 48402 50258 48414
rect 20414 48354 20466 48366
rect 20066 48302 20078 48354
rect 20130 48302 20142 48354
rect 20414 48290 20466 48302
rect 20638 48354 20690 48366
rect 20638 48290 20690 48302
rect 22094 48354 22146 48366
rect 22094 48290 22146 48302
rect 22318 48354 22370 48366
rect 22318 48290 22370 48302
rect 24558 48354 24610 48366
rect 24558 48290 24610 48302
rect 25566 48354 25618 48366
rect 25566 48290 25618 48302
rect 47070 48354 47122 48366
rect 47070 48290 47122 48302
rect 48750 48354 48802 48366
rect 48750 48290 48802 48302
rect 21310 48242 21362 48254
rect 21074 48190 21086 48242
rect 21138 48190 21150 48242
rect 21310 48178 21362 48190
rect 21646 48242 21698 48254
rect 23102 48242 23154 48254
rect 24446 48242 24498 48254
rect 25790 48242 25842 48254
rect 22642 48190 22654 48242
rect 22706 48190 22718 48242
rect 23986 48190 23998 48242
rect 24050 48190 24062 48242
rect 25218 48190 25230 48242
rect 25282 48190 25294 48242
rect 21646 48178 21698 48190
rect 23102 48178 23154 48190
rect 24446 48178 24498 48190
rect 25790 48178 25842 48190
rect 26238 48242 26290 48254
rect 26238 48178 26290 48190
rect 26462 48242 26514 48254
rect 26462 48178 26514 48190
rect 26910 48242 26962 48254
rect 26910 48178 26962 48190
rect 27582 48242 27634 48254
rect 40126 48242 40178 48254
rect 31938 48190 31950 48242
rect 32002 48190 32014 48242
rect 27582 48178 27634 48190
rect 40126 48178 40178 48190
rect 42478 48242 42530 48254
rect 46510 48242 46562 48254
rect 42914 48190 42926 48242
rect 42978 48190 42990 48242
rect 42478 48178 42530 48190
rect 46510 48178 46562 48190
rect 46846 48242 46898 48254
rect 46846 48178 46898 48190
rect 49870 48242 49922 48254
rect 51090 48190 51102 48242
rect 51154 48190 51166 48242
rect 49870 48178 49922 48190
rect 19518 48130 19570 48142
rect 21422 48130 21474 48142
rect 20738 48078 20750 48130
rect 20802 48078 20814 48130
rect 19518 48066 19570 48078
rect 21422 48066 21474 48078
rect 31614 48130 31666 48142
rect 31614 48066 31666 48078
rect 41022 48130 41074 48142
rect 41022 48066 41074 48078
rect 41806 48130 41858 48142
rect 46174 48130 46226 48142
rect 43586 48078 43598 48130
rect 43650 48078 43662 48130
rect 45714 48078 45726 48130
rect 45778 48078 45790 48130
rect 41806 48066 41858 48078
rect 46174 48066 46226 48078
rect 48190 48130 48242 48142
rect 48190 48066 48242 48078
rect 49310 48130 49362 48142
rect 49310 48066 49362 48078
rect 19742 48018 19794 48030
rect 19742 47954 19794 47966
rect 24222 48018 24274 48030
rect 24222 47954 24274 47966
rect 31950 48018 32002 48030
rect 31950 47954 32002 47966
rect 48974 48018 49026 48030
rect 48974 47954 49026 47966
rect 53006 48018 53058 48030
rect 53006 47954 53058 47966
rect 1344 47850 53648 47884
rect 1344 47798 4478 47850
rect 4530 47798 4582 47850
rect 4634 47798 4686 47850
rect 4738 47798 35198 47850
rect 35250 47798 35302 47850
rect 35354 47798 35406 47850
rect 35458 47798 53648 47850
rect 1344 47764 53648 47798
rect 43038 47682 43090 47694
rect 26562 47630 26574 47682
rect 26626 47630 26638 47682
rect 51314 47630 51326 47682
rect 51378 47679 51390 47682
rect 51538 47679 51550 47682
rect 51378 47633 51550 47679
rect 51378 47630 51390 47633
rect 51538 47630 51550 47633
rect 51602 47630 51614 47682
rect 43038 47618 43090 47630
rect 25342 47570 25394 47582
rect 38558 47570 38610 47582
rect 24098 47518 24110 47570
rect 24162 47518 24174 47570
rect 32050 47518 32062 47570
rect 32114 47518 32126 47570
rect 33170 47518 33182 47570
rect 33234 47518 33246 47570
rect 35298 47518 35310 47570
rect 35362 47518 35374 47570
rect 49634 47518 49646 47570
rect 49698 47518 49710 47570
rect 51090 47518 51102 47570
rect 51154 47518 51166 47570
rect 25342 47506 25394 47518
rect 38558 47506 38610 47518
rect 14030 47458 14082 47470
rect 14030 47394 14082 47406
rect 14590 47458 14642 47470
rect 14590 47394 14642 47406
rect 19294 47458 19346 47470
rect 25678 47458 25730 47470
rect 26350 47458 26402 47470
rect 19618 47406 19630 47458
rect 19682 47406 19694 47458
rect 25106 47406 25118 47458
rect 25170 47406 25182 47458
rect 26002 47406 26014 47458
rect 26066 47406 26078 47458
rect 19294 47394 19346 47406
rect 25678 47394 25730 47406
rect 26350 47394 26402 47406
rect 27022 47458 27074 47470
rect 27022 47394 27074 47406
rect 27134 47458 27186 47470
rect 27134 47394 27186 47406
rect 28254 47458 28306 47470
rect 29138 47406 29150 47458
rect 29202 47406 29214 47458
rect 32386 47406 32398 47458
rect 32450 47406 32462 47458
rect 41570 47406 41582 47458
rect 41634 47406 41646 47458
rect 49970 47406 49982 47458
rect 50034 47406 50046 47458
rect 28254 47394 28306 47406
rect 14142 47346 14194 47358
rect 14142 47282 14194 47294
rect 19406 47346 19458 47358
rect 19406 47282 19458 47294
rect 23774 47346 23826 47358
rect 24782 47346 24834 47358
rect 24434 47294 24446 47346
rect 24498 47294 24510 47346
rect 23774 47282 23826 47294
rect 24782 47282 24834 47294
rect 25454 47346 25506 47358
rect 25454 47282 25506 47294
rect 27246 47346 27298 47358
rect 27246 47282 27298 47294
rect 27694 47346 27746 47358
rect 27694 47282 27746 47294
rect 27918 47346 27970 47358
rect 27918 47282 27970 47294
rect 28142 47346 28194 47358
rect 41918 47346 41970 47358
rect 29922 47294 29934 47346
rect 29986 47294 29998 47346
rect 28142 47282 28194 47294
rect 41918 47282 41970 47294
rect 42254 47346 42306 47358
rect 42254 47282 42306 47294
rect 42702 47346 42754 47358
rect 42702 47282 42754 47294
rect 42926 47346 42978 47358
rect 42926 47282 42978 47294
rect 48750 47346 48802 47358
rect 48750 47282 48802 47294
rect 50430 47346 50482 47358
rect 50430 47282 50482 47294
rect 50766 47346 50818 47358
rect 50766 47282 50818 47294
rect 14254 47234 14306 47246
rect 23998 47234 24050 47246
rect 18834 47182 18846 47234
rect 18898 47182 18910 47234
rect 14254 47170 14306 47182
rect 23998 47170 24050 47182
rect 26238 47234 26290 47246
rect 26238 47170 26290 47182
rect 35758 47234 35810 47246
rect 35758 47170 35810 47182
rect 41806 47234 41858 47246
rect 41806 47170 41858 47182
rect 42030 47234 42082 47246
rect 42030 47170 42082 47182
rect 46174 47234 46226 47246
rect 46174 47170 46226 47182
rect 48862 47234 48914 47246
rect 48862 47170 48914 47182
rect 49086 47234 49138 47246
rect 49086 47170 49138 47182
rect 50990 47234 51042 47246
rect 50990 47170 51042 47182
rect 51662 47234 51714 47246
rect 51662 47170 51714 47182
rect 1344 47066 53648 47100
rect 1344 47014 19838 47066
rect 19890 47014 19942 47066
rect 19994 47014 20046 47066
rect 20098 47014 50558 47066
rect 50610 47014 50662 47066
rect 50714 47014 50766 47066
rect 50818 47014 53648 47066
rect 1344 46980 53648 47014
rect 13246 46898 13298 46910
rect 27470 46898 27522 46910
rect 14690 46846 14702 46898
rect 14754 46846 14766 46898
rect 21074 46846 21086 46898
rect 21138 46846 21150 46898
rect 13246 46834 13298 46846
rect 27470 46834 27522 46846
rect 27694 46898 27746 46910
rect 27694 46834 27746 46846
rect 32286 46898 32338 46910
rect 32286 46834 32338 46846
rect 38670 46898 38722 46910
rect 40002 46846 40014 46898
rect 40066 46846 40078 46898
rect 38670 46834 38722 46846
rect 12014 46786 12066 46798
rect 12014 46722 12066 46734
rect 12238 46786 12290 46798
rect 12238 46722 12290 46734
rect 14030 46786 14082 46798
rect 20414 46786 20466 46798
rect 23438 46786 23490 46798
rect 20066 46734 20078 46786
rect 20130 46734 20142 46786
rect 20962 46734 20974 46786
rect 21026 46734 21038 46786
rect 14030 46722 14082 46734
rect 20414 46722 20466 46734
rect 23438 46722 23490 46734
rect 27358 46786 27410 46798
rect 30258 46734 30270 46786
rect 30322 46734 30334 46786
rect 30930 46734 30942 46786
rect 30994 46734 31006 46786
rect 33506 46734 33518 46786
rect 33570 46734 33582 46786
rect 51090 46734 51102 46786
rect 51154 46734 51166 46786
rect 27358 46722 27410 46734
rect 12350 46674 12402 46686
rect 12350 46610 12402 46622
rect 13134 46674 13186 46686
rect 13134 46610 13186 46622
rect 13358 46674 13410 46686
rect 13358 46610 13410 46622
rect 13806 46674 13858 46686
rect 13806 46610 13858 46622
rect 14254 46674 14306 46686
rect 14254 46610 14306 46622
rect 14478 46674 14530 46686
rect 14478 46610 14530 46622
rect 14702 46674 14754 46686
rect 14702 46610 14754 46622
rect 15038 46674 15090 46686
rect 20302 46674 20354 46686
rect 18946 46622 18958 46674
rect 19010 46622 19022 46674
rect 19618 46622 19630 46674
rect 19682 46622 19694 46674
rect 15038 46610 15090 46622
rect 20302 46610 20354 46622
rect 22542 46674 22594 46686
rect 30158 46674 30210 46686
rect 38894 46674 38946 46686
rect 24658 46622 24670 46674
rect 24722 46622 24734 46674
rect 33730 46622 33742 46674
rect 33794 46622 33806 46674
rect 35522 46622 35534 46674
rect 35586 46622 35598 46674
rect 22542 46610 22594 46622
rect 30158 46610 30210 46622
rect 38894 46610 38946 46622
rect 39342 46674 39394 46686
rect 48190 46674 48242 46686
rect 40226 46622 40238 46674
rect 40290 46622 40302 46674
rect 47170 46622 47182 46674
rect 47234 46622 47246 46674
rect 39342 46610 39394 46622
rect 48190 46610 48242 46622
rect 48750 46674 48802 46686
rect 50306 46622 50318 46674
rect 50370 46622 50382 46674
rect 48750 46610 48802 46622
rect 11902 46562 11954 46574
rect 11902 46498 11954 46510
rect 12798 46562 12850 46574
rect 12798 46498 12850 46510
rect 15150 46562 15202 46574
rect 15150 46498 15202 46510
rect 29934 46562 29986 46574
rect 38782 46562 38834 46574
rect 36194 46510 36206 46562
rect 36258 46510 36270 46562
rect 38322 46510 38334 46562
rect 38386 46510 38398 46562
rect 29934 46498 29986 46510
rect 38782 46498 38834 46510
rect 39678 46562 39730 46574
rect 47742 46562 47794 46574
rect 44370 46510 44382 46562
rect 44434 46510 44446 46562
rect 46498 46510 46510 46562
rect 46562 46510 46574 46562
rect 39678 46498 39730 46510
rect 47742 46498 47794 46510
rect 49310 46562 49362 46574
rect 49310 46498 49362 46510
rect 49982 46562 50034 46574
rect 53218 46510 53230 46562
rect 53282 46510 53294 46562
rect 49982 46498 50034 46510
rect 1344 46282 53648 46316
rect 1344 46230 4478 46282
rect 4530 46230 4582 46282
rect 4634 46230 4686 46282
rect 4738 46230 35198 46282
rect 35250 46230 35302 46282
rect 35354 46230 35406 46282
rect 35458 46230 53648 46282
rect 1344 46196 53648 46230
rect 44158 46114 44210 46126
rect 18946 46062 18958 46114
rect 19010 46111 19022 46114
rect 19282 46111 19294 46114
rect 19010 46065 19294 46111
rect 19010 46062 19022 46065
rect 19282 46062 19294 46065
rect 19346 46062 19358 46114
rect 21858 46062 21870 46114
rect 21922 46062 21934 46114
rect 44158 46050 44210 46062
rect 37102 46002 37154 46014
rect 11554 45950 11566 46002
rect 11618 45950 11630 46002
rect 14242 45950 14254 46002
rect 14306 45950 14318 46002
rect 18722 45950 18734 46002
rect 18786 45950 18798 46002
rect 22530 45950 22542 46002
rect 22594 45950 22606 46002
rect 37102 45938 37154 45950
rect 38558 46002 38610 46014
rect 42354 45950 42366 46002
rect 42418 45950 42430 46002
rect 38558 45938 38610 45950
rect 12014 45890 12066 45902
rect 33966 45890 34018 45902
rect 37550 45890 37602 45902
rect 8754 45838 8766 45890
rect 8818 45838 8830 45890
rect 14018 45838 14030 45890
rect 14082 45838 14094 45890
rect 15026 45838 15038 45890
rect 15090 45838 15102 45890
rect 15922 45838 15934 45890
rect 15986 45838 15998 45890
rect 22418 45838 22430 45890
rect 22482 45838 22494 45890
rect 22642 45838 22654 45890
rect 22706 45838 22718 45890
rect 34290 45838 34302 45890
rect 34354 45838 34366 45890
rect 12014 45826 12066 45838
rect 33966 45826 34018 45838
rect 37550 45826 37602 45838
rect 38222 45890 38274 45902
rect 42030 45890 42082 45902
rect 39778 45838 39790 45890
rect 39842 45838 39854 45890
rect 38222 45826 38274 45838
rect 42030 45826 42082 45838
rect 43038 45890 43090 45902
rect 43038 45826 43090 45838
rect 43262 45890 43314 45902
rect 43262 45826 43314 45838
rect 43374 45890 43426 45902
rect 43374 45826 43426 45838
rect 36990 45778 37042 45790
rect 9426 45726 9438 45778
rect 9490 45726 9502 45778
rect 14466 45726 14478 45778
rect 14530 45726 14542 45778
rect 16594 45726 16606 45778
rect 16658 45726 16670 45778
rect 24322 45726 24334 45778
rect 24386 45726 24398 45778
rect 24994 45726 25006 45778
rect 25058 45726 25070 45778
rect 36990 45714 37042 45726
rect 37326 45778 37378 45790
rect 37326 45714 37378 45726
rect 37886 45778 37938 45790
rect 37886 45714 37938 45726
rect 37998 45778 38050 45790
rect 41806 45778 41858 45790
rect 39554 45726 39566 45778
rect 39618 45726 39630 45778
rect 40562 45726 40574 45778
rect 40626 45726 40638 45778
rect 37998 45714 38050 45726
rect 41806 45714 41858 45726
rect 42366 45778 42418 45790
rect 42366 45714 42418 45726
rect 43150 45778 43202 45790
rect 43150 45714 43202 45726
rect 43822 45778 43874 45790
rect 43822 45714 43874 45726
rect 49086 45778 49138 45790
rect 49086 45714 49138 45726
rect 12126 45666 12178 45678
rect 12126 45602 12178 45614
rect 12238 45666 12290 45678
rect 12238 45602 12290 45614
rect 12462 45666 12514 45678
rect 12462 45602 12514 45614
rect 13582 45666 13634 45678
rect 13582 45602 13634 45614
rect 19182 45666 19234 45678
rect 19182 45602 19234 45614
rect 23998 45666 24050 45678
rect 23998 45602 24050 45614
rect 24670 45666 24722 45678
rect 24670 45602 24722 45614
rect 25454 45666 25506 45678
rect 25454 45602 25506 45614
rect 34078 45666 34130 45678
rect 34078 45602 34130 45614
rect 40238 45666 40290 45678
rect 40238 45602 40290 45614
rect 42254 45666 42306 45678
rect 42254 45602 42306 45614
rect 42926 45666 42978 45678
rect 42926 45602 42978 45614
rect 44046 45666 44098 45678
rect 44046 45602 44098 45614
rect 49198 45666 49250 45678
rect 49198 45602 49250 45614
rect 1344 45498 53648 45532
rect 1344 45446 19838 45498
rect 19890 45446 19942 45498
rect 19994 45446 20046 45498
rect 20098 45446 50558 45498
rect 50610 45446 50662 45498
rect 50714 45446 50766 45498
rect 50818 45446 53648 45498
rect 1344 45412 53648 45446
rect 11566 45330 11618 45342
rect 22878 45330 22930 45342
rect 36542 45330 36594 45342
rect 12450 45278 12462 45330
rect 12514 45278 12526 45330
rect 23202 45278 23214 45330
rect 23266 45278 23278 45330
rect 11566 45266 11618 45278
rect 22878 45266 22930 45278
rect 36542 45266 36594 45278
rect 37326 45330 37378 45342
rect 41134 45330 41186 45342
rect 37986 45278 37998 45330
rect 38050 45278 38062 45330
rect 37326 45266 37378 45278
rect 41134 45266 41186 45278
rect 43150 45330 43202 45342
rect 43150 45266 43202 45278
rect 49982 45330 50034 45342
rect 49982 45266 50034 45278
rect 11790 45218 11842 45230
rect 11790 45154 11842 45166
rect 14254 45218 14306 45230
rect 14254 45154 14306 45166
rect 14366 45218 14418 45230
rect 14366 45154 14418 45166
rect 18062 45218 18114 45230
rect 18062 45154 18114 45166
rect 18622 45218 18674 45230
rect 18622 45154 18674 45166
rect 19070 45218 19122 45230
rect 19070 45154 19122 45166
rect 33406 45218 33458 45230
rect 33406 45154 33458 45166
rect 33630 45218 33682 45230
rect 42926 45218 42978 45230
rect 38322 45166 38334 45218
rect 38386 45166 38398 45218
rect 38882 45166 38894 45218
rect 38946 45166 38958 45218
rect 39442 45166 39454 45218
rect 39506 45166 39518 45218
rect 33630 45154 33682 45166
rect 42926 45154 42978 45166
rect 48190 45218 48242 45230
rect 48190 45154 48242 45166
rect 50094 45218 50146 45230
rect 50094 45154 50146 45166
rect 11342 45106 11394 45118
rect 11342 45042 11394 45054
rect 11566 45106 11618 45118
rect 18286 45106 18338 45118
rect 12226 45054 12238 45106
rect 12290 45054 12302 45106
rect 14018 45054 14030 45106
rect 14082 45054 14094 45106
rect 11566 45042 11618 45054
rect 18286 45042 18338 45054
rect 18958 45106 19010 45118
rect 26014 45106 26066 45118
rect 32286 45106 32338 45118
rect 35646 45106 35698 45118
rect 22642 45054 22654 45106
rect 22706 45054 22718 45106
rect 23426 45054 23438 45106
rect 23490 45054 23502 45106
rect 32050 45054 32062 45106
rect 32114 45054 32126 45106
rect 34626 45054 34638 45106
rect 34690 45054 34702 45106
rect 35410 45054 35422 45106
rect 35474 45054 35486 45106
rect 18958 45042 19010 45054
rect 26014 45042 26066 45054
rect 32286 45042 32338 45054
rect 35646 45042 35698 45054
rect 35758 45106 35810 45118
rect 35758 45042 35810 45054
rect 37102 45106 37154 45118
rect 37102 45042 37154 45054
rect 37438 45106 37490 45118
rect 41358 45106 41410 45118
rect 38434 45054 38446 45106
rect 38498 45054 38510 45106
rect 38770 45054 38782 45106
rect 38834 45054 38846 45106
rect 40898 45054 40910 45106
rect 40962 45054 40974 45106
rect 37438 45042 37490 45054
rect 41358 45042 41410 45054
rect 41470 45106 41522 45118
rect 48974 45106 49026 45118
rect 49758 45106 49810 45118
rect 43810 45054 43822 45106
rect 43874 45054 43886 45106
rect 47842 45054 47854 45106
rect 47906 45054 47918 45106
rect 49186 45054 49198 45106
rect 49250 45054 49262 45106
rect 51090 45054 51102 45106
rect 51154 45054 51166 45106
rect 41470 45042 41522 45054
rect 48974 45042 49026 45054
rect 49758 45042 49810 45054
rect 15374 44994 15426 45006
rect 15374 44930 15426 44942
rect 18174 44994 18226 45006
rect 18174 44930 18226 44942
rect 19742 44994 19794 45006
rect 19742 44930 19794 44942
rect 24558 44994 24610 45006
rect 24558 44930 24610 44942
rect 31502 44994 31554 45006
rect 31502 44930 31554 44942
rect 34190 44994 34242 45006
rect 34190 44930 34242 44942
rect 41246 44994 41298 45006
rect 47070 44994 47122 45006
rect 43250 44942 43262 44994
rect 43314 44942 43326 44994
rect 44482 44942 44494 44994
rect 44546 44942 44558 44994
rect 46610 44942 46622 44994
rect 46674 44942 46686 44994
rect 41246 44930 41298 44942
rect 47070 44930 47122 44942
rect 47518 44994 47570 45006
rect 47518 44930 47570 44942
rect 48078 44994 48130 45006
rect 48078 44930 48130 44942
rect 48750 44994 48802 45006
rect 48750 44930 48802 44942
rect 19070 44882 19122 44894
rect 14802 44830 14814 44882
rect 14866 44830 14878 44882
rect 19070 44818 19122 44830
rect 26126 44882 26178 44894
rect 26126 44818 26178 44830
rect 33294 44882 33346 44894
rect 36206 44882 36258 44894
rect 34290 44830 34302 44882
rect 34354 44830 34366 44882
rect 33294 44818 33346 44830
rect 36206 44818 36258 44830
rect 36430 44882 36482 44894
rect 36430 44818 36482 44830
rect 53006 44882 53058 44894
rect 53006 44818 53058 44830
rect 1344 44714 53648 44748
rect 1344 44662 4478 44714
rect 4530 44662 4582 44714
rect 4634 44662 4686 44714
rect 4738 44662 35198 44714
rect 35250 44662 35302 44714
rect 35354 44662 35406 44714
rect 35458 44662 53648 44714
rect 1344 44628 53648 44662
rect 17278 44546 17330 44558
rect 17278 44482 17330 44494
rect 17614 44546 17666 44558
rect 17614 44482 17666 44494
rect 22094 44546 22146 44558
rect 22094 44482 22146 44494
rect 26910 44546 26962 44558
rect 26910 44482 26962 44494
rect 17726 44434 17778 44446
rect 17726 44370 17778 44382
rect 18622 44434 18674 44446
rect 18622 44370 18674 44382
rect 19406 44434 19458 44446
rect 19406 44370 19458 44382
rect 26126 44434 26178 44446
rect 32510 44434 32562 44446
rect 32050 44382 32062 44434
rect 32114 44382 32126 44434
rect 26126 44370 26178 44382
rect 32510 44370 32562 44382
rect 32846 44434 32898 44446
rect 32846 44370 32898 44382
rect 33966 44434 34018 44446
rect 48514 44382 48526 44434
rect 48578 44382 48590 44434
rect 33966 44370 34018 44382
rect 16830 44322 16882 44334
rect 16146 44270 16158 44322
rect 16210 44270 16222 44322
rect 16830 44258 16882 44270
rect 17390 44322 17442 44334
rect 17390 44258 17442 44270
rect 18174 44322 18226 44334
rect 18174 44258 18226 44270
rect 18846 44322 18898 44334
rect 18846 44258 18898 44270
rect 19854 44322 19906 44334
rect 19854 44258 19906 44270
rect 20078 44322 20130 44334
rect 20078 44258 20130 44270
rect 22206 44322 22258 44334
rect 22206 44258 22258 44270
rect 22878 44322 22930 44334
rect 25454 44322 25506 44334
rect 23426 44270 23438 44322
rect 23490 44270 23502 44322
rect 22878 44258 22930 44270
rect 25454 44258 25506 44270
rect 25790 44322 25842 44334
rect 29138 44270 29150 44322
rect 29202 44270 29214 44322
rect 34738 44270 34750 44322
rect 34802 44270 34814 44322
rect 35746 44270 35758 44322
rect 35810 44270 35822 44322
rect 48962 44270 48974 44322
rect 49026 44270 49038 44322
rect 25790 44258 25842 44270
rect 18398 44210 18450 44222
rect 25118 44210 25170 44222
rect 49422 44210 49474 44222
rect 16370 44158 16382 44210
rect 16434 44158 16446 44210
rect 22530 44158 22542 44210
rect 22594 44158 22606 44210
rect 29922 44158 29934 44210
rect 29986 44158 29998 44210
rect 34850 44158 34862 44210
rect 34914 44158 34926 44210
rect 36418 44158 36430 44210
rect 36482 44158 36494 44210
rect 18398 44146 18450 44158
rect 25118 44146 25170 44158
rect 49422 44146 49474 44158
rect 50542 44210 50594 44222
rect 50542 44146 50594 44158
rect 11566 44098 11618 44110
rect 11566 44034 11618 44046
rect 19518 44098 19570 44110
rect 19518 44034 19570 44046
rect 19966 44098 20018 44110
rect 19966 44034 20018 44046
rect 20302 44098 20354 44110
rect 20302 44034 20354 44046
rect 22094 44098 22146 44110
rect 25454 44098 25506 44110
rect 23202 44046 23214 44098
rect 23266 44046 23278 44098
rect 22094 44034 22146 44046
rect 25454 44034 25506 44046
rect 26014 44098 26066 44110
rect 26014 44034 26066 44046
rect 26238 44098 26290 44110
rect 26238 44034 26290 44046
rect 26462 44098 26514 44110
rect 26462 44034 26514 44046
rect 27022 44098 27074 44110
rect 27022 44034 27074 44046
rect 27134 44098 27186 44110
rect 27134 44034 27186 44046
rect 32958 44098 33010 44110
rect 32958 44034 33010 44046
rect 33406 44098 33458 44110
rect 38670 44098 38722 44110
rect 36306 44046 36318 44098
rect 36370 44046 36382 44098
rect 33406 44034 33458 44046
rect 38670 44034 38722 44046
rect 49982 44098 50034 44110
rect 49982 44034 50034 44046
rect 50878 44098 50930 44110
rect 50878 44034 50930 44046
rect 1344 43930 53648 43964
rect 1344 43878 19838 43930
rect 19890 43878 19942 43930
rect 19994 43878 20046 43930
rect 20098 43878 50558 43930
rect 50610 43878 50662 43930
rect 50714 43878 50766 43930
rect 50818 43878 53648 43930
rect 1344 43844 53648 43878
rect 18062 43762 18114 43774
rect 11218 43710 11230 43762
rect 11282 43710 11294 43762
rect 18062 43698 18114 43710
rect 20190 43762 20242 43774
rect 26126 43762 26178 43774
rect 21410 43710 21422 43762
rect 21474 43710 21486 43762
rect 20190 43698 20242 43710
rect 26126 43698 26178 43710
rect 29374 43762 29426 43774
rect 38894 43762 38946 43774
rect 33730 43710 33742 43762
rect 33794 43710 33806 43762
rect 34402 43710 34414 43762
rect 34466 43710 34478 43762
rect 29374 43698 29426 43710
rect 38894 43698 38946 43710
rect 46062 43762 46114 43774
rect 46062 43698 46114 43710
rect 11790 43650 11842 43662
rect 11790 43586 11842 43598
rect 12350 43650 12402 43662
rect 12350 43586 12402 43598
rect 12574 43650 12626 43662
rect 12574 43586 12626 43598
rect 14030 43650 14082 43662
rect 14030 43586 14082 43598
rect 14142 43650 14194 43662
rect 14142 43586 14194 43598
rect 18734 43650 18786 43662
rect 18734 43586 18786 43598
rect 20078 43650 20130 43662
rect 20078 43586 20130 43598
rect 20750 43650 20802 43662
rect 20750 43586 20802 43598
rect 21086 43650 21138 43662
rect 21086 43586 21138 43598
rect 26798 43650 26850 43662
rect 26798 43586 26850 43598
rect 27918 43650 27970 43662
rect 28578 43598 28590 43650
rect 28642 43598 28654 43650
rect 49634 43598 49646 43650
rect 49698 43598 49710 43650
rect 51090 43598 51102 43650
rect 51154 43598 51166 43650
rect 27918 43586 27970 43598
rect 10894 43538 10946 43550
rect 10894 43474 10946 43486
rect 11566 43538 11618 43550
rect 11566 43474 11618 43486
rect 12238 43538 12290 43550
rect 12238 43474 12290 43486
rect 12686 43538 12738 43550
rect 14702 43538 14754 43550
rect 14354 43486 14366 43538
rect 14418 43486 14430 43538
rect 12686 43474 12738 43486
rect 14702 43474 14754 43486
rect 18286 43538 18338 43550
rect 18286 43474 18338 43486
rect 18958 43538 19010 43550
rect 18958 43474 19010 43486
rect 20414 43538 20466 43550
rect 20414 43474 20466 43486
rect 25566 43538 25618 43550
rect 27134 43538 27186 43550
rect 25890 43486 25902 43538
rect 25954 43486 25966 43538
rect 25566 43474 25618 43486
rect 27134 43474 27186 43486
rect 27358 43538 27410 43550
rect 29262 43538 29314 43550
rect 34078 43538 34130 43550
rect 28354 43486 28366 43538
rect 28418 43486 28430 43538
rect 33506 43486 33518 43538
rect 33570 43486 33582 43538
rect 27358 43474 27410 43486
rect 29262 43474 29314 43486
rect 34078 43474 34130 43486
rect 38782 43538 38834 43550
rect 38782 43474 38834 43486
rect 39118 43538 39170 43550
rect 39118 43474 39170 43486
rect 45950 43538 46002 43550
rect 45950 43474 46002 43486
rect 46286 43538 46338 43550
rect 46286 43474 46338 43486
rect 49086 43538 49138 43550
rect 49086 43474 49138 43486
rect 49310 43538 49362 43550
rect 50306 43486 50318 43538
rect 50370 43486 50382 43538
rect 49310 43474 49362 43486
rect 12014 43426 12066 43438
rect 12014 43362 12066 43374
rect 18510 43426 18562 43438
rect 18510 43362 18562 43374
rect 19854 43426 19906 43438
rect 19854 43362 19906 43374
rect 25790 43426 25842 43438
rect 25790 43362 25842 43374
rect 27246 43426 27298 43438
rect 27246 43362 27298 43374
rect 34862 43426 34914 43438
rect 34862 43362 34914 43374
rect 48302 43426 48354 43438
rect 53218 43374 53230 43426
rect 53282 43374 53294 43426
rect 48302 43362 48354 43374
rect 29038 43314 29090 43326
rect 29038 43250 29090 43262
rect 29374 43314 29426 43326
rect 29374 43250 29426 43262
rect 1344 43146 53648 43180
rect 1344 43094 4478 43146
rect 4530 43094 4582 43146
rect 4634 43094 4686 43146
rect 4738 43094 35198 43146
rect 35250 43094 35302 43146
rect 35354 43094 35406 43146
rect 35458 43094 53648 43146
rect 1344 43060 53648 43094
rect 14030 42978 14082 42990
rect 14030 42914 14082 42926
rect 14366 42978 14418 42990
rect 29710 42978 29762 42990
rect 15250 42926 15262 42978
rect 15314 42926 15326 42978
rect 14366 42914 14418 42926
rect 29710 42914 29762 42926
rect 33966 42978 34018 42990
rect 33966 42914 34018 42926
rect 38670 42978 38722 42990
rect 38670 42914 38722 42926
rect 12238 42866 12290 42878
rect 9650 42814 9662 42866
rect 9714 42814 9726 42866
rect 11778 42814 11790 42866
rect 11842 42814 11854 42866
rect 12238 42802 12290 42814
rect 16046 42866 16098 42878
rect 23650 42814 23662 42866
rect 23714 42814 23726 42866
rect 43138 42814 43150 42866
rect 43202 42814 43214 42866
rect 16046 42802 16098 42814
rect 14702 42754 14754 42766
rect 24110 42754 24162 42766
rect 8866 42702 8878 42754
rect 8930 42702 8942 42754
rect 15362 42702 15374 42754
rect 15426 42702 15438 42754
rect 14702 42690 14754 42702
rect 24110 42690 24162 42702
rect 33070 42754 33122 42766
rect 33070 42690 33122 42702
rect 33294 42754 33346 42766
rect 33294 42690 33346 42702
rect 33518 42754 33570 42766
rect 33518 42690 33570 42702
rect 36990 42754 37042 42766
rect 36990 42690 37042 42702
rect 37774 42754 37826 42766
rect 37774 42690 37826 42702
rect 38446 42754 38498 42766
rect 44270 42754 44322 42766
rect 40338 42702 40350 42754
rect 40402 42702 40414 42754
rect 38446 42690 38498 42702
rect 44270 42690 44322 42702
rect 44830 42754 44882 42766
rect 44830 42690 44882 42702
rect 45390 42754 45442 42766
rect 45390 42690 45442 42702
rect 13806 42642 13858 42654
rect 37102 42642 37154 42654
rect 14914 42590 14926 42642
rect 14978 42590 14990 42642
rect 13806 42578 13858 42590
rect 37102 42578 37154 42590
rect 37662 42642 37714 42654
rect 39678 42642 39730 42654
rect 43486 42642 43538 42654
rect 38994 42590 39006 42642
rect 39058 42590 39070 42642
rect 39330 42590 39342 42642
rect 39394 42590 39406 42642
rect 41010 42590 41022 42642
rect 41074 42590 41086 42642
rect 37662 42578 37714 42590
rect 39678 42578 39730 42590
rect 43486 42578 43538 42590
rect 45502 42642 45554 42654
rect 45502 42578 45554 42590
rect 23550 42530 23602 42542
rect 15138 42478 15150 42530
rect 15202 42478 15214 42530
rect 23550 42466 23602 42478
rect 23774 42530 23826 42542
rect 23774 42466 23826 42478
rect 28590 42530 28642 42542
rect 28590 42466 28642 42478
rect 29822 42530 29874 42542
rect 29822 42466 29874 42478
rect 29934 42530 29986 42542
rect 29934 42466 29986 42478
rect 30494 42530 30546 42542
rect 30494 42466 30546 42478
rect 32286 42530 32338 42542
rect 32286 42466 32338 42478
rect 32734 42530 32786 42542
rect 32734 42466 32786 42478
rect 37326 42530 37378 42542
rect 37326 42466 37378 42478
rect 37438 42530 37490 42542
rect 37438 42466 37490 42478
rect 43822 42530 43874 42542
rect 43822 42466 43874 42478
rect 44942 42530 44994 42542
rect 44942 42466 44994 42478
rect 45166 42530 45218 42542
rect 45166 42466 45218 42478
rect 45726 42530 45778 42542
rect 45726 42466 45778 42478
rect 49982 42530 50034 42542
rect 49982 42466 50034 42478
rect 1344 42362 53648 42396
rect 1344 42310 19838 42362
rect 19890 42310 19942 42362
rect 19994 42310 20046 42362
rect 20098 42310 50558 42362
rect 50610 42310 50662 42362
rect 50714 42310 50766 42362
rect 50818 42310 53648 42362
rect 1344 42276 53648 42310
rect 12686 42194 12738 42206
rect 12686 42130 12738 42142
rect 14142 42194 14194 42206
rect 14142 42130 14194 42142
rect 14366 42194 14418 42206
rect 14366 42130 14418 42142
rect 15038 42194 15090 42206
rect 15038 42130 15090 42142
rect 23550 42194 23602 42206
rect 33182 42194 33234 42206
rect 27010 42142 27022 42194
rect 27074 42142 27086 42194
rect 23550 42130 23602 42142
rect 33182 42130 33234 42142
rect 38446 42194 38498 42206
rect 38446 42130 38498 42142
rect 40014 42194 40066 42206
rect 40014 42130 40066 42142
rect 41134 42194 41186 42206
rect 41134 42130 41186 42142
rect 43262 42194 43314 42206
rect 43262 42130 43314 42142
rect 49870 42194 49922 42206
rect 49870 42130 49922 42142
rect 14590 42082 14642 42094
rect 14590 42018 14642 42030
rect 15150 42082 15202 42094
rect 38334 42082 38386 42094
rect 29810 42030 29822 42082
rect 29874 42030 29886 42082
rect 15150 42018 15202 42030
rect 38334 42018 38386 42030
rect 39902 42082 39954 42094
rect 39902 42018 39954 42030
rect 43374 42082 43426 42094
rect 43374 42018 43426 42030
rect 12350 41970 12402 41982
rect 5058 41918 5070 41970
rect 5122 41918 5134 41970
rect 12350 41906 12402 41918
rect 22990 41970 23042 41982
rect 23774 41970 23826 41982
rect 23314 41918 23326 41970
rect 23378 41918 23390 41970
rect 22990 41906 23042 41918
rect 23774 41906 23826 41918
rect 23886 41970 23938 41982
rect 23886 41906 23938 41918
rect 26126 41970 26178 41982
rect 26126 41906 26178 41918
rect 26350 41970 26402 41982
rect 26350 41906 26402 41918
rect 26798 41970 26850 41982
rect 26798 41906 26850 41918
rect 27358 41970 27410 41982
rect 33518 41970 33570 41982
rect 29138 41918 29150 41970
rect 29202 41918 29214 41970
rect 27358 41906 27410 41918
rect 33518 41906 33570 41918
rect 38670 41970 38722 41982
rect 38670 41906 38722 41918
rect 40238 41970 40290 41982
rect 41246 41970 41298 41982
rect 48862 41970 48914 41982
rect 40898 41918 40910 41970
rect 40962 41918 40974 41970
rect 48066 41918 48078 41970
rect 48130 41918 48142 41970
rect 40238 41906 40290 41918
rect 41246 41906 41298 41918
rect 48862 41906 48914 41918
rect 49310 41970 49362 41982
rect 50418 41918 50430 41970
rect 50482 41918 50494 41970
rect 49310 41906 49362 41918
rect 8318 41858 8370 41870
rect 5730 41806 5742 41858
rect 5794 41806 5806 41858
rect 7858 41806 7870 41858
rect 7922 41806 7934 41858
rect 8318 41794 8370 41806
rect 23662 41858 23714 41870
rect 23662 41794 23714 41806
rect 24446 41858 24498 41870
rect 24446 41794 24498 41806
rect 26574 41858 26626 41870
rect 26574 41794 26626 41806
rect 31950 41858 32002 41870
rect 31950 41794 32002 41806
rect 36654 41858 36706 41870
rect 45266 41806 45278 41858
rect 45330 41806 45342 41858
rect 47394 41806 47406 41858
rect 47458 41806 47470 41858
rect 49858 41806 49870 41858
rect 49922 41806 49934 41858
rect 51090 41806 51102 41858
rect 51154 41806 51166 41858
rect 53218 41806 53230 41858
rect 53282 41806 53294 41858
rect 36654 41794 36706 41806
rect 14478 41746 14530 41758
rect 14478 41682 14530 41694
rect 15038 41746 15090 41758
rect 24334 41746 24386 41758
rect 22642 41694 22654 41746
rect 22706 41743 22718 41746
rect 23090 41743 23102 41746
rect 22706 41697 23102 41743
rect 22706 41694 22718 41697
rect 23090 41694 23102 41697
rect 23154 41694 23166 41746
rect 15038 41682 15090 41694
rect 24334 41682 24386 41694
rect 33182 41746 33234 41758
rect 33182 41682 33234 41694
rect 33294 41746 33346 41758
rect 33294 41682 33346 41694
rect 43262 41746 43314 41758
rect 43262 41682 43314 41694
rect 49646 41746 49698 41758
rect 49646 41682 49698 41694
rect 1344 41578 53648 41612
rect 1344 41526 4478 41578
rect 4530 41526 4582 41578
rect 4634 41526 4686 41578
rect 4738 41526 35198 41578
rect 35250 41526 35302 41578
rect 35354 41526 35406 41578
rect 35458 41526 53648 41578
rect 1344 41492 53648 41526
rect 14814 41410 14866 41422
rect 14814 41346 14866 41358
rect 26462 41410 26514 41422
rect 26462 41346 26514 41358
rect 26798 41410 26850 41422
rect 26798 41346 26850 41358
rect 32398 41298 32450 41310
rect 49086 41298 49138 41310
rect 17042 41246 17054 41298
rect 17106 41246 17118 41298
rect 19170 41246 19182 41298
rect 19234 41246 19246 41298
rect 24770 41246 24782 41298
rect 24834 41246 24846 41298
rect 36418 41246 36430 41298
rect 36482 41246 36494 41298
rect 32398 41234 32450 41246
rect 49086 41234 49138 41246
rect 51886 41298 51938 41310
rect 51886 41234 51938 41246
rect 14366 41186 14418 41198
rect 14366 41122 14418 41134
rect 14702 41186 14754 41198
rect 26574 41186 26626 41198
rect 37326 41186 37378 41198
rect 15138 41134 15150 41186
rect 15202 41134 15214 41186
rect 16370 41134 16382 41186
rect 16434 41134 16446 41186
rect 22194 41134 22206 41186
rect 22258 41134 22270 41186
rect 22754 41134 22766 41186
rect 22818 41134 22830 41186
rect 26002 41134 26014 41186
rect 26066 41134 26078 41186
rect 33506 41134 33518 41186
rect 33570 41134 33582 41186
rect 14702 41122 14754 41134
rect 26574 41122 26626 41134
rect 37326 41122 37378 41134
rect 45614 41186 45666 41198
rect 45614 41122 45666 41134
rect 48526 41186 48578 41198
rect 48526 41122 48578 41134
rect 49198 41186 49250 41198
rect 49970 41134 49982 41186
rect 50034 41134 50046 41186
rect 49198 41122 49250 41134
rect 36990 41074 37042 41086
rect 23426 41022 23438 41074
rect 23490 41022 23502 41074
rect 24546 41022 24558 41074
rect 24610 41022 24622 41074
rect 34290 41022 34302 41074
rect 34354 41022 34366 41074
rect 36990 41010 37042 41022
rect 37102 41074 37154 41086
rect 37102 41010 37154 41022
rect 37550 41074 37602 41086
rect 37550 41010 37602 41022
rect 45278 41074 45330 41086
rect 45278 41010 45330 41022
rect 45838 41074 45890 41086
rect 45838 41010 45890 41022
rect 14478 40962 14530 40974
rect 14478 40898 14530 40910
rect 15598 40962 15650 40974
rect 15598 40898 15650 40910
rect 19630 40962 19682 40974
rect 26462 40962 26514 40974
rect 22418 40910 22430 40962
rect 22482 40910 22494 40962
rect 19630 40898 19682 40910
rect 26462 40898 26514 40910
rect 27358 40962 27410 40974
rect 27358 40898 27410 40910
rect 40574 40962 40626 40974
rect 40574 40898 40626 40910
rect 41806 40962 41858 40974
rect 41806 40898 41858 40910
rect 45726 40962 45778 40974
rect 45726 40898 45778 40910
rect 48414 40962 48466 40974
rect 48414 40898 48466 40910
rect 48974 40962 49026 40974
rect 48974 40898 49026 40910
rect 1344 40794 53648 40828
rect 1344 40742 19838 40794
rect 19890 40742 19942 40794
rect 19994 40742 20046 40794
rect 20098 40742 50558 40794
rect 50610 40742 50662 40794
rect 50714 40742 50766 40794
rect 50818 40742 53648 40794
rect 1344 40708 53648 40742
rect 5742 40626 5794 40638
rect 5742 40562 5794 40574
rect 15374 40626 15426 40638
rect 15374 40562 15426 40574
rect 22654 40626 22706 40638
rect 24334 40626 24386 40638
rect 23314 40574 23326 40626
rect 23378 40574 23390 40626
rect 22654 40562 22706 40574
rect 24334 40562 24386 40574
rect 38894 40626 38946 40638
rect 38894 40562 38946 40574
rect 42030 40626 42082 40638
rect 42030 40562 42082 40574
rect 44046 40626 44098 40638
rect 44046 40562 44098 40574
rect 44270 40626 44322 40638
rect 44270 40562 44322 40574
rect 7982 40514 8034 40526
rect 22990 40514 23042 40526
rect 19730 40462 19742 40514
rect 19794 40462 19806 40514
rect 7982 40450 8034 40462
rect 22990 40450 23042 40462
rect 23886 40514 23938 40526
rect 23886 40450 23938 40462
rect 24222 40514 24274 40526
rect 35310 40514 35362 40526
rect 40126 40514 40178 40526
rect 26562 40462 26574 40514
rect 26626 40462 26638 40514
rect 38546 40462 38558 40514
rect 38610 40462 38622 40514
rect 24222 40450 24274 40462
rect 35310 40450 35362 40462
rect 40126 40450 40178 40462
rect 41470 40514 41522 40526
rect 43710 40514 43762 40526
rect 42354 40462 42366 40514
rect 42418 40462 42430 40514
rect 41470 40450 41522 40462
rect 43710 40450 43762 40462
rect 5406 40402 5458 40414
rect 5406 40338 5458 40350
rect 5742 40402 5794 40414
rect 5742 40338 5794 40350
rect 5966 40402 6018 40414
rect 5966 40338 6018 40350
rect 8318 40402 8370 40414
rect 8318 40338 8370 40350
rect 16606 40402 16658 40414
rect 16606 40338 16658 40350
rect 18622 40402 18674 40414
rect 23326 40402 23378 40414
rect 19058 40350 19070 40402
rect 19122 40350 19134 40402
rect 18622 40338 18674 40350
rect 23326 40338 23378 40350
rect 23438 40402 23490 40414
rect 23438 40338 23490 40350
rect 23662 40402 23714 40414
rect 23662 40338 23714 40350
rect 24558 40402 24610 40414
rect 29150 40402 29202 40414
rect 33294 40402 33346 40414
rect 40014 40402 40066 40414
rect 25890 40350 25902 40402
rect 25954 40350 25966 40402
rect 31938 40350 31950 40402
rect 32002 40350 32014 40402
rect 32162 40350 32174 40402
rect 32226 40350 32238 40402
rect 38098 40350 38110 40402
rect 38162 40350 38174 40402
rect 24558 40338 24610 40350
rect 29150 40338 29202 40350
rect 33294 40338 33346 40350
rect 40014 40338 40066 40350
rect 40798 40402 40850 40414
rect 40798 40338 40850 40350
rect 41134 40402 41186 40414
rect 41134 40338 41186 40350
rect 43934 40402 43986 40414
rect 44482 40350 44494 40402
rect 44546 40350 44558 40402
rect 50642 40350 50654 40402
rect 50706 40350 50718 40402
rect 43934 40338 43986 40350
rect 15486 40290 15538 40302
rect 32398 40290 32450 40302
rect 41022 40290 41074 40302
rect 21858 40238 21870 40290
rect 21922 40238 21934 40290
rect 28690 40238 28702 40290
rect 28754 40238 28766 40290
rect 35746 40238 35758 40290
rect 35810 40238 35822 40290
rect 46834 40238 46846 40290
rect 46898 40238 46910 40290
rect 15486 40226 15538 40238
rect 32398 40226 32450 40238
rect 41022 40226 41074 40238
rect 40126 40178 40178 40190
rect 40126 40114 40178 40126
rect 53006 40178 53058 40190
rect 53006 40114 53058 40126
rect 1344 40010 53648 40044
rect 1344 39958 4478 40010
rect 4530 39958 4582 40010
rect 4634 39958 4686 40010
rect 4738 39958 35198 40010
rect 35250 39958 35302 40010
rect 35354 39958 35406 40010
rect 35458 39958 53648 40010
rect 1344 39924 53648 39958
rect 5966 39842 6018 39854
rect 5966 39778 6018 39790
rect 6526 39842 6578 39854
rect 6526 39778 6578 39790
rect 8430 39842 8482 39854
rect 8430 39778 8482 39790
rect 37102 39842 37154 39854
rect 37102 39778 37154 39790
rect 23998 39730 24050 39742
rect 12786 39678 12798 39730
rect 12850 39678 12862 39730
rect 14242 39678 14254 39730
rect 14306 39678 14318 39730
rect 16370 39678 16382 39730
rect 16434 39678 16446 39730
rect 17378 39678 17390 39730
rect 17442 39678 17454 39730
rect 23998 39666 24050 39678
rect 27918 39730 27970 39742
rect 38434 39678 38446 39730
rect 38498 39678 38510 39730
rect 40562 39678 40574 39730
rect 40626 39678 40638 39730
rect 46722 39678 46734 39730
rect 46786 39678 46798 39730
rect 27918 39666 27970 39678
rect 9326 39618 9378 39630
rect 9326 39554 9378 39566
rect 9550 39618 9602 39630
rect 19294 39618 19346 39630
rect 41806 39618 41858 39630
rect 9874 39566 9886 39618
rect 9938 39566 9950 39618
rect 13570 39566 13582 39618
rect 13634 39566 13646 39618
rect 17042 39566 17054 39618
rect 17106 39566 17118 39618
rect 18946 39566 18958 39618
rect 19010 39566 19022 39618
rect 28354 39566 28366 39618
rect 28418 39566 28430 39618
rect 41346 39566 41358 39618
rect 41410 39566 41422 39618
rect 9550 39554 9602 39566
rect 19294 39554 19346 39566
rect 41806 39554 41858 39566
rect 44046 39618 44098 39630
rect 44046 39554 44098 39566
rect 44718 39618 44770 39630
rect 44718 39554 44770 39566
rect 45166 39618 45218 39630
rect 50318 39618 50370 39630
rect 49634 39566 49646 39618
rect 49698 39566 49710 39618
rect 45166 39554 45218 39566
rect 50318 39554 50370 39566
rect 50766 39618 50818 39630
rect 50766 39554 50818 39566
rect 50878 39618 50930 39630
rect 50878 39554 50930 39566
rect 51326 39618 51378 39630
rect 51326 39554 51378 39566
rect 4958 39506 5010 39518
rect 4958 39442 5010 39454
rect 5630 39506 5682 39518
rect 5630 39442 5682 39454
rect 6078 39506 6130 39518
rect 6078 39442 6130 39454
rect 6414 39506 6466 39518
rect 6414 39442 6466 39454
rect 6526 39506 6578 39518
rect 6526 39442 6578 39454
rect 8094 39506 8146 39518
rect 8094 39442 8146 39454
rect 8542 39506 8594 39518
rect 8542 39442 8594 39454
rect 8990 39506 9042 39518
rect 8990 39442 9042 39454
rect 9438 39506 9490 39518
rect 17726 39506 17778 39518
rect 10658 39454 10670 39506
rect 10722 39454 10734 39506
rect 9438 39442 9490 39454
rect 17726 39442 17778 39454
rect 19406 39506 19458 39518
rect 19406 39442 19458 39454
rect 36206 39506 36258 39518
rect 36206 39442 36258 39454
rect 37102 39506 37154 39518
rect 37102 39442 37154 39454
rect 37214 39506 37266 39518
rect 37214 39442 37266 39454
rect 45390 39506 45442 39518
rect 45390 39442 45442 39454
rect 46062 39506 46114 39518
rect 52110 39506 52162 39518
rect 48850 39454 48862 39506
rect 48914 39454 48926 39506
rect 46062 39442 46114 39454
rect 52110 39442 52162 39454
rect 5070 39394 5122 39406
rect 5070 39330 5122 39342
rect 5854 39394 5906 39406
rect 5854 39330 5906 39342
rect 8318 39394 8370 39406
rect 8318 39330 8370 39342
rect 36318 39394 36370 39406
rect 36318 39330 36370 39342
rect 36542 39394 36594 39406
rect 36542 39330 36594 39342
rect 44158 39394 44210 39406
rect 44158 39330 44210 39342
rect 44382 39394 44434 39406
rect 44382 39330 44434 39342
rect 44942 39394 44994 39406
rect 44942 39330 44994 39342
rect 46174 39394 46226 39406
rect 46174 39330 46226 39342
rect 46398 39394 46450 39406
rect 46398 39330 46450 39342
rect 50206 39394 50258 39406
rect 50206 39330 50258 39342
rect 50990 39394 51042 39406
rect 50990 39330 51042 39342
rect 51438 39394 51490 39406
rect 51438 39330 51490 39342
rect 51550 39394 51602 39406
rect 51550 39330 51602 39342
rect 1344 39226 53648 39260
rect 1344 39174 19838 39226
rect 19890 39174 19942 39226
rect 19994 39174 20046 39226
rect 20098 39174 50558 39226
rect 50610 39174 50662 39226
rect 50714 39174 50766 39226
rect 50818 39174 53648 39226
rect 1344 39140 53648 39174
rect 7198 39058 7250 39070
rect 7198 38994 7250 39006
rect 9886 39058 9938 39070
rect 9886 38994 9938 39006
rect 10110 39058 10162 39070
rect 10110 38994 10162 39006
rect 13022 39058 13074 39070
rect 13022 38994 13074 39006
rect 19518 39058 19570 39070
rect 19518 38994 19570 39006
rect 34862 39058 34914 39070
rect 34862 38994 34914 39006
rect 46398 39058 46450 39070
rect 46398 38994 46450 39006
rect 46958 39058 47010 39070
rect 46958 38994 47010 39006
rect 7982 38946 8034 38958
rect 7982 38882 8034 38894
rect 8094 38946 8146 38958
rect 8094 38882 8146 38894
rect 19742 38946 19794 38958
rect 47070 38946 47122 38958
rect 22306 38894 22318 38946
rect 22370 38894 22382 38946
rect 30930 38894 30942 38946
rect 30994 38894 31006 38946
rect 32386 38894 32398 38946
rect 32450 38894 32462 38946
rect 44930 38894 44942 38946
rect 44994 38894 45006 38946
rect 19742 38882 19794 38894
rect 47070 38882 47122 38894
rect 47294 38946 47346 38958
rect 51090 38894 51102 38946
rect 51154 38894 51166 38946
rect 47294 38882 47346 38894
rect 7534 38834 7586 38846
rect 7534 38770 7586 38782
rect 8206 38834 8258 38846
rect 8206 38770 8258 38782
rect 9774 38834 9826 38846
rect 17950 38834 18002 38846
rect 16370 38782 16382 38834
rect 16434 38782 16446 38834
rect 16594 38782 16606 38834
rect 16658 38782 16670 38834
rect 9774 38770 9826 38782
rect 17950 38770 18002 38782
rect 19854 38834 19906 38846
rect 30494 38834 30546 38846
rect 33294 38834 33346 38846
rect 46622 38834 46674 38846
rect 20850 38782 20862 38834
rect 20914 38782 20926 38834
rect 21634 38782 21646 38834
rect 21698 38782 21710 38834
rect 30034 38782 30046 38834
rect 30098 38782 30110 38834
rect 30818 38782 30830 38834
rect 30882 38782 30894 38834
rect 32498 38782 32510 38834
rect 32562 38782 32574 38834
rect 33730 38782 33742 38834
rect 33794 38782 33806 38834
rect 37762 38782 37774 38834
rect 37826 38782 37838 38834
rect 45714 38782 45726 38834
rect 45778 38782 45790 38834
rect 50418 38782 50430 38834
rect 50482 38782 50494 38834
rect 19854 38770 19906 38782
rect 30494 38770 30546 38782
rect 33294 38770 33346 38782
rect 46622 38770 46674 38782
rect 16830 38722 16882 38734
rect 17614 38722 17666 38734
rect 17378 38670 17390 38722
rect 17442 38719 17454 38722
rect 17442 38673 17551 38719
rect 17442 38670 17454 38673
rect 16830 38658 16882 38670
rect 8642 38558 8654 38610
rect 8706 38558 8718 38610
rect 17505 38607 17551 38673
rect 17614 38658 17666 38670
rect 20190 38722 20242 38734
rect 24446 38722 24498 38734
rect 21074 38670 21086 38722
rect 21138 38670 21150 38722
rect 20190 38658 20242 38670
rect 24446 38658 24498 38670
rect 29262 38722 29314 38734
rect 29586 38670 29598 38722
rect 29650 38670 29662 38722
rect 32050 38670 32062 38722
rect 32114 38670 32126 38722
rect 33618 38670 33630 38722
rect 33682 38670 33694 38722
rect 36306 38670 36318 38722
rect 36370 38670 36382 38722
rect 42802 38670 42814 38722
rect 42866 38670 42878 38722
rect 53218 38670 53230 38722
rect 53282 38670 53294 38722
rect 29262 38658 29314 38670
rect 17938 38607 17950 38610
rect 17505 38561 17950 38607
rect 17938 38558 17950 38561
rect 18002 38558 18014 38610
rect 1344 38442 53648 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 53648 38442
rect 1344 38356 53648 38390
rect 5966 38274 6018 38286
rect 5966 38210 6018 38222
rect 8766 38274 8818 38286
rect 8766 38210 8818 38222
rect 17950 38274 18002 38286
rect 17950 38210 18002 38222
rect 31390 38162 31442 38174
rect 44270 38162 44322 38174
rect 8530 38110 8542 38162
rect 8594 38110 8606 38162
rect 19954 38110 19966 38162
rect 20018 38110 20030 38162
rect 36418 38110 36430 38162
rect 36482 38110 36494 38162
rect 45938 38110 45950 38162
rect 46002 38110 46014 38162
rect 31390 38098 31442 38110
rect 44270 38098 44322 38110
rect 6078 38050 6130 38062
rect 6078 37986 6130 37998
rect 18062 38050 18114 38062
rect 18062 37986 18114 37998
rect 18286 38050 18338 38062
rect 18286 37986 18338 37998
rect 18510 38050 18562 38062
rect 18510 37986 18562 37998
rect 18622 38050 18674 38062
rect 20190 38050 20242 38062
rect 26350 38050 26402 38062
rect 28478 38050 28530 38062
rect 19618 37998 19630 38050
rect 19682 37998 19694 38050
rect 25778 37998 25790 38050
rect 25842 37998 25854 38050
rect 28130 37998 28142 38050
rect 28194 37998 28206 38050
rect 18622 37986 18674 37998
rect 20190 37986 20242 37998
rect 26350 37986 26402 37998
rect 28478 37986 28530 37998
rect 30046 38050 30098 38062
rect 30046 37986 30098 37998
rect 30494 38050 30546 38062
rect 32286 38050 32338 38062
rect 36990 38050 37042 38062
rect 30706 37998 30718 38050
rect 30770 37998 30782 38050
rect 33618 37998 33630 38050
rect 33682 37998 33694 38050
rect 30494 37986 30546 37998
rect 32286 37986 32338 37998
rect 36990 37986 37042 37998
rect 37326 38050 37378 38062
rect 37326 37986 37378 37998
rect 37550 38050 37602 38062
rect 44818 37998 44830 38050
rect 44882 37998 44894 38050
rect 37550 37986 37602 37998
rect 4958 37938 5010 37950
rect 4958 37874 5010 37886
rect 5070 37938 5122 37950
rect 5070 37874 5122 37886
rect 5966 37938 6018 37950
rect 5966 37874 6018 37886
rect 9550 37938 9602 37950
rect 9550 37874 9602 37886
rect 9662 37938 9714 37950
rect 26462 37938 26514 37950
rect 19058 37886 19070 37938
rect 19122 37886 19134 37938
rect 20626 37886 20638 37938
rect 20690 37886 20702 37938
rect 9662 37874 9714 37886
rect 26462 37874 26514 37886
rect 28590 37938 28642 37950
rect 28590 37874 28642 37886
rect 31950 37938 32002 37950
rect 31950 37874 32002 37886
rect 32062 37938 32114 37950
rect 37102 37938 37154 37950
rect 34290 37886 34302 37938
rect 34354 37886 34366 37938
rect 32062 37874 32114 37886
rect 37102 37874 37154 37886
rect 38894 37938 38946 37950
rect 40898 37886 40910 37938
rect 40962 37886 40974 37938
rect 38894 37874 38946 37886
rect 4734 37826 4786 37838
rect 4734 37762 4786 37774
rect 8542 37826 8594 37838
rect 8542 37762 8594 37774
rect 9886 37826 9938 37838
rect 9886 37762 9938 37774
rect 21422 37826 21474 37838
rect 21422 37762 21474 37774
rect 26910 37826 26962 37838
rect 26910 37762 26962 37774
rect 29262 37826 29314 37838
rect 29262 37762 29314 37774
rect 32958 37826 33010 37838
rect 32958 37762 33010 37774
rect 37998 37826 38050 37838
rect 37998 37762 38050 37774
rect 38558 37826 38610 37838
rect 38558 37762 38610 37774
rect 38782 37826 38834 37838
rect 38782 37762 38834 37774
rect 41246 37826 41298 37838
rect 41246 37762 41298 37774
rect 1344 37658 53648 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 50558 37658
rect 50610 37606 50662 37658
rect 50714 37606 50766 37658
rect 50818 37606 53648 37658
rect 1344 37572 53648 37606
rect 5854 37490 5906 37502
rect 5854 37426 5906 37438
rect 5966 37490 6018 37502
rect 8878 37490 8930 37502
rect 7522 37438 7534 37490
rect 7586 37438 7598 37490
rect 5966 37426 6018 37438
rect 8878 37426 8930 37438
rect 8990 37490 9042 37502
rect 49310 37490 49362 37502
rect 29362 37438 29374 37490
rect 29426 37438 29438 37490
rect 8990 37426 9042 37438
rect 49310 37426 49362 37438
rect 5294 37378 5346 37390
rect 5294 37314 5346 37326
rect 5518 37378 5570 37390
rect 5518 37314 5570 37326
rect 9550 37378 9602 37390
rect 9550 37314 9602 37326
rect 9662 37378 9714 37390
rect 9662 37314 9714 37326
rect 9886 37378 9938 37390
rect 9886 37314 9938 37326
rect 10446 37378 10498 37390
rect 10446 37314 10498 37326
rect 15934 37378 15986 37390
rect 15934 37314 15986 37326
rect 18510 37378 18562 37390
rect 18510 37314 18562 37326
rect 26798 37378 26850 37390
rect 43262 37378 43314 37390
rect 28018 37326 28030 37378
rect 28082 37326 28094 37378
rect 29474 37326 29486 37378
rect 29538 37326 29550 37378
rect 26798 37314 26850 37326
rect 43262 37314 43314 37326
rect 43822 37378 43874 37390
rect 43822 37314 43874 37326
rect 44046 37378 44098 37390
rect 44046 37314 44098 37326
rect 44158 37378 44210 37390
rect 44158 37314 44210 37326
rect 49086 37378 49138 37390
rect 49086 37314 49138 37326
rect 4846 37266 4898 37278
rect 1810 37214 1822 37266
rect 1874 37214 1886 37266
rect 4846 37202 4898 37214
rect 6078 37266 6130 37278
rect 6078 37202 6130 37214
rect 6526 37266 6578 37278
rect 6526 37202 6578 37214
rect 8318 37266 8370 37278
rect 8318 37202 8370 37214
rect 8766 37266 8818 37278
rect 8766 37202 8818 37214
rect 9998 37266 10050 37278
rect 9998 37202 10050 37214
rect 10222 37266 10274 37278
rect 10222 37202 10274 37214
rect 10670 37266 10722 37278
rect 15822 37266 15874 37278
rect 10994 37214 11006 37266
rect 11058 37214 11070 37266
rect 11778 37214 11790 37266
rect 11842 37214 11854 37266
rect 15250 37214 15262 37266
rect 15314 37214 15326 37266
rect 10670 37202 10722 37214
rect 15822 37202 15874 37214
rect 16494 37266 16546 37278
rect 26238 37266 26290 37278
rect 43150 37266 43202 37278
rect 19058 37214 19070 37266
rect 19122 37214 19134 37266
rect 25554 37214 25566 37266
rect 25618 37214 25630 37266
rect 28466 37214 28478 37266
rect 28530 37214 28542 37266
rect 28914 37214 28926 37266
rect 28978 37214 28990 37266
rect 37538 37214 37550 37266
rect 37602 37214 37614 37266
rect 16494 37202 16546 37214
rect 26238 37202 26290 37214
rect 43150 37202 43202 37214
rect 43710 37266 43762 37278
rect 43710 37202 43762 37214
rect 48638 37266 48690 37278
rect 50418 37214 50430 37266
rect 50482 37214 50494 37266
rect 48638 37202 48690 37214
rect 5070 37154 5122 37166
rect 2482 37102 2494 37154
rect 2546 37102 2558 37154
rect 4610 37102 4622 37154
rect 4674 37102 4686 37154
rect 5070 37090 5122 37102
rect 6974 37154 7026 37166
rect 14366 37154 14418 37166
rect 20078 37154 20130 37166
rect 36430 37154 36482 37166
rect 13906 37102 13918 37154
rect 13970 37102 13982 37154
rect 19394 37102 19406 37154
rect 19458 37102 19470 37154
rect 25330 37102 25342 37154
rect 25394 37102 25406 37154
rect 6974 37090 7026 37102
rect 14366 37090 14418 37102
rect 20078 37090 20130 37102
rect 36430 37090 36482 37102
rect 37102 37154 37154 37166
rect 42702 37154 42754 37166
rect 38210 37102 38222 37154
rect 38274 37102 38286 37154
rect 40338 37102 40350 37154
rect 40402 37102 40414 37154
rect 37102 37090 37154 37102
rect 42702 37090 42754 37102
rect 43486 37154 43538 37166
rect 43486 37090 43538 37102
rect 48190 37154 48242 37166
rect 48190 37090 48242 37102
rect 49198 37154 49250 37166
rect 51090 37102 51102 37154
rect 51154 37102 51166 37154
rect 53218 37102 53230 37154
rect 53282 37102 53294 37154
rect 49198 37090 49250 37102
rect 7198 37042 7250 37054
rect 7198 36978 7250 36990
rect 1344 36874 53648 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 53648 36874
rect 1344 36788 53648 36822
rect 5742 36706 5794 36718
rect 5742 36642 5794 36654
rect 9438 36706 9490 36718
rect 9438 36642 9490 36654
rect 18398 36594 18450 36606
rect 5954 36542 5966 36594
rect 6018 36542 6030 36594
rect 18398 36530 18450 36542
rect 18734 36594 18786 36606
rect 18734 36530 18786 36542
rect 28590 36594 28642 36606
rect 28590 36530 28642 36542
rect 38894 36594 38946 36606
rect 51214 36594 51266 36606
rect 48962 36542 48974 36594
rect 49026 36542 49038 36594
rect 38894 36530 38946 36542
rect 51214 36530 51266 36542
rect 15486 36482 15538 36494
rect 18846 36482 18898 36494
rect 38670 36482 38722 36494
rect 6066 36430 6078 36482
rect 6130 36430 6142 36482
rect 9426 36430 9438 36482
rect 9490 36430 9502 36482
rect 15138 36430 15150 36482
rect 15202 36430 15214 36482
rect 17714 36430 17726 36482
rect 17778 36430 17790 36482
rect 18162 36430 18174 36482
rect 18226 36430 18238 36482
rect 19170 36430 19182 36482
rect 19234 36430 19246 36482
rect 21634 36430 21646 36482
rect 21698 36430 21710 36482
rect 28130 36430 28142 36482
rect 28194 36430 28206 36482
rect 28354 36430 28366 36482
rect 28418 36430 28430 36482
rect 30258 36430 30270 36482
rect 30322 36430 30334 36482
rect 15486 36418 15538 36430
rect 18846 36418 18898 36430
rect 38670 36418 38722 36430
rect 39118 36482 39170 36494
rect 50094 36482 50146 36494
rect 46162 36430 46174 36482
rect 46226 36430 46238 36482
rect 39118 36418 39170 36430
rect 50094 36418 50146 36430
rect 50542 36482 50594 36494
rect 50542 36418 50594 36430
rect 50766 36482 50818 36494
rect 50766 36418 50818 36430
rect 9102 36370 9154 36382
rect 9102 36306 9154 36318
rect 15598 36370 15650 36382
rect 15598 36306 15650 36318
rect 16046 36370 16098 36382
rect 36206 36370 36258 36382
rect 22418 36318 22430 36370
rect 22482 36318 22494 36370
rect 30930 36318 30942 36370
rect 30994 36318 31006 36370
rect 16046 36306 16098 36318
rect 36206 36306 36258 36318
rect 39342 36370 39394 36382
rect 50654 36370 50706 36382
rect 46834 36318 46846 36370
rect 46898 36318 46910 36370
rect 39342 36306 39394 36318
rect 50654 36306 50706 36318
rect 51102 36370 51154 36382
rect 51102 36306 51154 36318
rect 4846 36258 4898 36270
rect 4846 36194 4898 36206
rect 10894 36258 10946 36270
rect 10894 36194 10946 36206
rect 20190 36258 20242 36270
rect 29262 36258 29314 36270
rect 33742 36258 33794 36270
rect 24658 36206 24670 36258
rect 24722 36206 24734 36258
rect 33170 36206 33182 36258
rect 33234 36206 33246 36258
rect 20190 36194 20242 36206
rect 29262 36194 29314 36206
rect 33742 36194 33794 36206
rect 35758 36258 35810 36270
rect 35758 36194 35810 36206
rect 37214 36258 37266 36270
rect 37214 36194 37266 36206
rect 39790 36258 39842 36270
rect 39790 36194 39842 36206
rect 51326 36258 51378 36270
rect 51326 36194 51378 36206
rect 1344 36090 53648 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 50558 36090
rect 50610 36038 50662 36090
rect 50714 36038 50766 36090
rect 50818 36038 53648 36090
rect 1344 36004 53648 36038
rect 4846 35922 4898 35934
rect 21870 35922 21922 35934
rect 7522 35870 7534 35922
rect 7586 35870 7598 35922
rect 4846 35858 4898 35870
rect 21870 35858 21922 35870
rect 22318 35922 22370 35934
rect 22318 35858 22370 35870
rect 22878 35922 22930 35934
rect 22878 35858 22930 35870
rect 38894 35922 38946 35934
rect 38894 35858 38946 35870
rect 46286 35922 46338 35934
rect 46286 35858 46338 35870
rect 5518 35810 5570 35822
rect 5518 35746 5570 35758
rect 8318 35810 8370 35822
rect 8318 35746 8370 35758
rect 8430 35810 8482 35822
rect 8430 35746 8482 35758
rect 22542 35810 22594 35822
rect 46622 35810 46674 35822
rect 36530 35758 36542 35810
rect 36594 35758 36606 35810
rect 38434 35758 38446 35810
rect 38498 35758 38510 35810
rect 44482 35758 44494 35810
rect 44546 35758 44558 35810
rect 49746 35758 49758 35810
rect 49810 35758 49822 35810
rect 22542 35746 22594 35758
rect 46622 35746 46674 35758
rect 5630 35698 5682 35710
rect 5630 35634 5682 35646
rect 7870 35698 7922 35710
rect 7870 35634 7922 35646
rect 8542 35698 8594 35710
rect 22206 35698 22258 35710
rect 16258 35646 16270 35698
rect 16322 35646 16334 35698
rect 8542 35634 8594 35646
rect 22206 35634 22258 35646
rect 22654 35698 22706 35710
rect 22654 35634 22706 35646
rect 23102 35698 23154 35710
rect 23102 35634 23154 35646
rect 23326 35698 23378 35710
rect 45950 35698 46002 35710
rect 33058 35646 33070 35698
rect 33122 35646 33134 35698
rect 36866 35646 36878 35698
rect 36930 35646 36942 35698
rect 37314 35646 37326 35698
rect 37378 35646 37390 35698
rect 37874 35646 37886 35698
rect 37938 35646 37950 35698
rect 38210 35646 38222 35698
rect 38274 35646 38286 35698
rect 45266 35646 45278 35698
rect 45330 35646 45342 35698
rect 23326 35634 23378 35646
rect 45950 35634 46002 35646
rect 46286 35698 46338 35710
rect 46286 35634 46338 35646
rect 49422 35698 49474 35710
rect 50642 35646 50654 35698
rect 50706 35646 50718 35698
rect 49422 35634 49474 35646
rect 15822 35586 15874 35598
rect 23774 35586 23826 35598
rect 35982 35586 36034 35598
rect 16594 35534 16606 35586
rect 16658 35534 16670 35586
rect 33842 35534 33854 35586
rect 33906 35534 33918 35586
rect 15822 35522 15874 35534
rect 23774 35522 23826 35534
rect 35982 35522 36034 35534
rect 41582 35586 41634 35598
rect 49086 35586 49138 35598
rect 42354 35534 42366 35586
rect 42418 35534 42430 35586
rect 41582 35522 41634 35534
rect 49086 35522 49138 35534
rect 5518 35474 5570 35486
rect 53006 35474 53058 35486
rect 8978 35422 8990 35474
rect 9042 35422 9054 35474
rect 5518 35410 5570 35422
rect 53006 35410 53058 35422
rect 1344 35306 53648 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 53648 35306
rect 1344 35220 53648 35254
rect 32734 35026 32786 35038
rect 4610 34974 4622 35026
rect 4674 34974 4686 35026
rect 28354 34974 28366 35026
rect 28418 34974 28430 35026
rect 32162 34974 32174 35026
rect 32226 34974 32238 35026
rect 32734 34962 32786 34974
rect 5518 34914 5570 34926
rect 1810 34862 1822 34914
rect 1874 34862 1886 34914
rect 5518 34850 5570 34862
rect 5854 34914 5906 34926
rect 5854 34850 5906 34862
rect 6190 34914 6242 34926
rect 18846 34914 18898 34926
rect 8754 34862 8766 34914
rect 8818 34862 8830 34914
rect 14354 34862 14366 34914
rect 14418 34862 14430 34914
rect 14802 34862 14814 34914
rect 14866 34862 14878 34914
rect 18498 34862 18510 34914
rect 18562 34862 18574 34914
rect 6190 34850 6242 34862
rect 18846 34850 18898 34862
rect 24558 34914 24610 34926
rect 36206 34914 36258 34926
rect 25330 34862 25342 34914
rect 25394 34862 25406 34914
rect 29250 34862 29262 34914
rect 29314 34862 29326 34914
rect 24558 34850 24610 34862
rect 36206 34850 36258 34862
rect 37886 34914 37938 34926
rect 40014 34914 40066 34926
rect 38322 34862 38334 34914
rect 38386 34862 38398 34914
rect 39106 34862 39118 34914
rect 39170 34862 39182 34914
rect 37886 34850 37938 34862
rect 40014 34850 40066 34862
rect 40574 34914 40626 34926
rect 40574 34850 40626 34862
rect 41582 34914 41634 34926
rect 41582 34850 41634 34862
rect 43934 34914 43986 34926
rect 43934 34850 43986 34862
rect 44830 34914 44882 34926
rect 44830 34850 44882 34862
rect 5070 34802 5122 34814
rect 2482 34750 2494 34802
rect 2546 34750 2558 34802
rect 5070 34738 5122 34750
rect 5742 34802 5794 34814
rect 9886 34802 9938 34814
rect 8978 34750 8990 34802
rect 9042 34750 9054 34802
rect 9538 34750 9550 34802
rect 9602 34750 9614 34802
rect 5742 34738 5794 34750
rect 9886 34738 9938 34750
rect 15038 34802 15090 34814
rect 15038 34738 15090 34750
rect 18958 34802 19010 34814
rect 42590 34802 42642 34814
rect 26114 34750 26126 34802
rect 26178 34750 26190 34802
rect 29922 34750 29934 34802
rect 29986 34750 29998 34802
rect 37314 34750 37326 34802
rect 37378 34750 37390 34802
rect 39330 34750 39342 34802
rect 39394 34750 39406 34802
rect 18958 34738 19010 34750
rect 42590 34738 42642 34750
rect 42702 34802 42754 34814
rect 42702 34738 42754 34750
rect 43822 34802 43874 34814
rect 43822 34738 43874 34750
rect 44942 34802 44994 34814
rect 44942 34738 44994 34750
rect 4958 34690 5010 34702
rect 4958 34626 5010 34638
rect 8094 34690 8146 34702
rect 8094 34626 8146 34638
rect 15486 34690 15538 34702
rect 15486 34626 15538 34638
rect 19406 34690 19458 34702
rect 19406 34626 19458 34638
rect 24222 34690 24274 34702
rect 24222 34626 24274 34638
rect 24670 34690 24722 34702
rect 24670 34626 24722 34638
rect 24894 34690 24946 34702
rect 24894 34626 24946 34638
rect 35758 34690 35810 34702
rect 35758 34626 35810 34638
rect 37102 34690 37154 34702
rect 41246 34690 41298 34702
rect 42366 34690 42418 34702
rect 39442 34638 39454 34690
rect 39506 34638 39518 34690
rect 40898 34638 40910 34690
rect 40962 34638 40974 34690
rect 41906 34638 41918 34690
rect 41970 34638 41982 34690
rect 37102 34626 37154 34638
rect 41246 34626 41298 34638
rect 42366 34626 42418 34638
rect 43598 34690 43650 34702
rect 43598 34626 43650 34638
rect 45166 34690 45218 34702
rect 45166 34626 45218 34638
rect 1344 34522 53648 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 50558 34522
rect 50610 34470 50662 34522
rect 50714 34470 50766 34522
rect 50818 34470 53648 34522
rect 1344 34436 53648 34470
rect 4958 34354 5010 34366
rect 4958 34290 5010 34302
rect 5182 34354 5234 34366
rect 5182 34290 5234 34302
rect 5966 34354 6018 34366
rect 5966 34290 6018 34302
rect 25790 34354 25842 34366
rect 25790 34290 25842 34302
rect 28702 34354 28754 34366
rect 28702 34290 28754 34302
rect 38670 34354 38722 34366
rect 38670 34290 38722 34302
rect 39790 34354 39842 34366
rect 39790 34290 39842 34302
rect 43822 34354 43874 34366
rect 43822 34290 43874 34302
rect 49086 34354 49138 34366
rect 49086 34290 49138 34302
rect 49310 34354 49362 34366
rect 49310 34290 49362 34302
rect 18734 34242 18786 34254
rect 18734 34178 18786 34190
rect 30382 34242 30434 34254
rect 49758 34242 49810 34254
rect 42130 34190 42142 34242
rect 42194 34190 42206 34242
rect 30382 34178 30434 34190
rect 49758 34178 49810 34190
rect 5518 34130 5570 34142
rect 5518 34066 5570 34078
rect 5854 34130 5906 34142
rect 5854 34066 5906 34078
rect 6078 34130 6130 34142
rect 6078 34066 6130 34078
rect 6526 34130 6578 34142
rect 13806 34130 13858 34142
rect 10546 34078 10558 34130
rect 10610 34078 10622 34130
rect 6526 34066 6578 34078
rect 13806 34066 13858 34078
rect 15486 34130 15538 34142
rect 25454 34130 25506 34142
rect 20514 34078 20526 34130
rect 20578 34078 20590 34130
rect 15486 34066 15538 34078
rect 25454 34066 25506 34078
rect 25902 34130 25954 34142
rect 25902 34066 25954 34078
rect 26014 34130 26066 34142
rect 26014 34066 26066 34078
rect 30270 34130 30322 34142
rect 30270 34066 30322 34078
rect 30606 34130 30658 34142
rect 38894 34130 38946 34142
rect 38434 34078 38446 34130
rect 38498 34078 38510 34130
rect 30606 34066 30658 34078
rect 38894 34066 38946 34078
rect 39006 34130 39058 34142
rect 39006 34066 39058 34078
rect 39902 34130 39954 34142
rect 42478 34130 42530 34142
rect 41010 34078 41022 34130
rect 41074 34078 41086 34130
rect 39902 34066 39954 34078
rect 42478 34066 42530 34078
rect 42814 34130 42866 34142
rect 42814 34066 42866 34078
rect 43374 34130 43426 34142
rect 43374 34066 43426 34078
rect 43710 34130 43762 34142
rect 45378 34078 45390 34130
rect 45442 34078 45454 34130
rect 48738 34078 48750 34130
rect 48802 34078 48814 34130
rect 50306 34078 50318 34130
rect 50370 34078 50382 34130
rect 43710 34066 43762 34078
rect 5294 34018 5346 34030
rect 18286 34018 18338 34030
rect 11218 33966 11230 34018
rect 11282 33966 11294 34018
rect 13346 33966 13358 34018
rect 13410 33966 13422 34018
rect 5294 33954 5346 33966
rect 18286 33954 18338 33966
rect 19182 34018 19234 34030
rect 24670 34018 24722 34030
rect 21186 33966 21198 34018
rect 21250 33966 21262 34018
rect 23314 33966 23326 34018
rect 23378 33966 23390 34018
rect 19182 33954 19234 33966
rect 24670 33954 24722 33966
rect 30942 34018 30994 34030
rect 30942 33954 30994 33966
rect 36654 34018 36706 34030
rect 36654 33954 36706 33966
rect 38110 34018 38162 34030
rect 38110 33954 38162 33966
rect 38782 34018 38834 34030
rect 49198 34018 49250 34030
rect 41346 33966 41358 34018
rect 41410 33966 41422 34018
rect 46050 33966 46062 34018
rect 46114 33966 46126 34018
rect 48178 33966 48190 34018
rect 48242 33966 48254 34018
rect 38782 33954 38834 33966
rect 49198 33954 49250 33966
rect 49870 34018 49922 34030
rect 51090 33966 51102 34018
rect 51154 33966 51166 34018
rect 53218 33966 53230 34018
rect 53282 33966 53294 34018
rect 49870 33954 49922 33966
rect 39790 33906 39842 33918
rect 39790 33842 39842 33854
rect 43822 33906 43874 33918
rect 43822 33842 43874 33854
rect 49982 33906 50034 33918
rect 49982 33842 50034 33854
rect 1344 33738 53648 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 53648 33738
rect 1344 33652 53648 33686
rect 9214 33570 9266 33582
rect 9214 33506 9266 33518
rect 29598 33570 29650 33582
rect 29598 33506 29650 33518
rect 30158 33570 30210 33582
rect 30158 33506 30210 33518
rect 33182 33570 33234 33582
rect 33182 33506 33234 33518
rect 11678 33458 11730 33470
rect 21422 33458 21474 33470
rect 41694 33458 41746 33470
rect 9538 33406 9550 33458
rect 9602 33406 9614 33458
rect 16706 33406 16718 33458
rect 16770 33406 16782 33458
rect 31042 33406 31054 33458
rect 31106 33406 31118 33458
rect 11678 33394 11730 33406
rect 21422 33394 21474 33406
rect 41694 33394 41746 33406
rect 45502 33458 45554 33470
rect 45502 33394 45554 33406
rect 48414 33458 48466 33470
rect 48414 33394 48466 33406
rect 50430 33458 50482 33470
rect 50430 33394 50482 33406
rect 5742 33346 5794 33358
rect 6302 33346 6354 33358
rect 5954 33294 5966 33346
rect 6018 33294 6030 33346
rect 5742 33282 5794 33294
rect 6302 33282 6354 33294
rect 10446 33346 10498 33358
rect 10446 33282 10498 33294
rect 10894 33346 10946 33358
rect 19406 33346 19458 33358
rect 14690 33294 14702 33346
rect 14754 33294 14766 33346
rect 15026 33294 15038 33346
rect 15090 33294 15102 33346
rect 17938 33294 17950 33346
rect 18002 33294 18014 33346
rect 18834 33294 18846 33346
rect 18898 33294 18910 33346
rect 10894 33282 10946 33294
rect 19406 33282 19458 33294
rect 19966 33346 20018 33358
rect 19966 33282 20018 33294
rect 20862 33346 20914 33358
rect 20862 33282 20914 33294
rect 21198 33346 21250 33358
rect 21198 33282 21250 33294
rect 23214 33346 23266 33358
rect 23214 33282 23266 33294
rect 25902 33346 25954 33358
rect 25902 33282 25954 33294
rect 29710 33346 29762 33358
rect 29710 33282 29762 33294
rect 29934 33346 29986 33358
rect 29934 33282 29986 33294
rect 30718 33346 30770 33358
rect 30718 33282 30770 33294
rect 33854 33346 33906 33358
rect 33854 33282 33906 33294
rect 45614 33346 45666 33358
rect 45614 33282 45666 33294
rect 45950 33346 46002 33358
rect 45950 33282 46002 33294
rect 49870 33346 49922 33358
rect 49870 33282 49922 33294
rect 50542 33346 50594 33358
rect 50542 33282 50594 33294
rect 5630 33234 5682 33246
rect 5630 33170 5682 33182
rect 10110 33234 10162 33246
rect 10110 33170 10162 33182
rect 10670 33234 10722 33246
rect 10670 33170 10722 33182
rect 11230 33234 11282 33246
rect 11230 33170 11282 33182
rect 15262 33234 15314 33246
rect 15262 33170 15314 33182
rect 19518 33234 19570 33246
rect 19518 33170 19570 33182
rect 20526 33234 20578 33246
rect 20526 33170 20578 33182
rect 21646 33234 21698 33246
rect 21646 33170 21698 33182
rect 21870 33234 21922 33246
rect 21870 33170 21922 33182
rect 23550 33234 23602 33246
rect 23550 33170 23602 33182
rect 25566 33234 25618 33246
rect 25566 33170 25618 33182
rect 33294 33234 33346 33246
rect 33294 33170 33346 33182
rect 33518 33234 33570 33246
rect 33518 33170 33570 33182
rect 33742 33234 33794 33246
rect 33742 33170 33794 33182
rect 34302 33234 34354 33246
rect 34302 33170 34354 33182
rect 45390 33234 45442 33246
rect 45390 33170 45442 33182
rect 6414 33122 6466 33134
rect 6414 33058 6466 33070
rect 6638 33122 6690 33134
rect 8318 33122 8370 33134
rect 7970 33070 7982 33122
rect 8034 33070 8046 33122
rect 6638 33058 6690 33070
rect 8318 33058 8370 33070
rect 8766 33122 8818 33134
rect 8766 33058 8818 33070
rect 9438 33122 9490 33134
rect 9438 33058 9490 33070
rect 10222 33122 10274 33134
rect 10222 33058 10274 33070
rect 10894 33122 10946 33134
rect 10894 33058 10946 33070
rect 20638 33122 20690 33134
rect 20638 33058 20690 33070
rect 23438 33122 23490 33134
rect 23438 33058 23490 33070
rect 24110 33122 24162 33134
rect 24110 33058 24162 33070
rect 25678 33122 25730 33134
rect 25678 33058 25730 33070
rect 26350 33122 26402 33134
rect 26350 33058 26402 33070
rect 29598 33122 29650 33134
rect 29598 33058 29650 33070
rect 30270 33122 30322 33134
rect 30270 33058 30322 33070
rect 30494 33122 30546 33134
rect 30494 33058 30546 33070
rect 31054 33122 31106 33134
rect 31054 33058 31106 33070
rect 31278 33122 31330 33134
rect 31278 33058 31330 33070
rect 32846 33122 32898 33134
rect 32846 33058 32898 33070
rect 33070 33122 33122 33134
rect 33070 33058 33122 33070
rect 40686 33122 40738 33134
rect 40686 33058 40738 33070
rect 50318 33122 50370 33134
rect 50318 33058 50370 33070
rect 1344 32954 53648 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 50558 32954
rect 50610 32902 50662 32954
rect 50714 32902 50766 32954
rect 50818 32902 53648 32954
rect 1344 32868 53648 32902
rect 9886 32786 9938 32798
rect 22766 32786 22818 32798
rect 19058 32734 19070 32786
rect 19122 32734 19134 32786
rect 20850 32734 20862 32786
rect 20914 32734 20926 32786
rect 9886 32722 9938 32734
rect 22766 32722 22818 32734
rect 26238 32786 26290 32798
rect 26238 32722 26290 32734
rect 31166 32786 31218 32798
rect 34078 32786 34130 32798
rect 33394 32734 33406 32786
rect 33458 32734 33470 32786
rect 31166 32722 31218 32734
rect 34078 32722 34130 32734
rect 41246 32786 41298 32798
rect 41246 32722 41298 32734
rect 43374 32786 43426 32798
rect 43586 32734 43598 32786
rect 43650 32734 43662 32786
rect 43374 32722 43426 32734
rect 5294 32674 5346 32686
rect 5294 32610 5346 32622
rect 5630 32674 5682 32686
rect 5630 32610 5682 32622
rect 6078 32674 6130 32686
rect 6078 32610 6130 32622
rect 6190 32674 6242 32686
rect 6190 32610 6242 32622
rect 6414 32674 6466 32686
rect 6414 32610 6466 32622
rect 6638 32674 6690 32686
rect 6638 32610 6690 32622
rect 9550 32674 9602 32686
rect 9550 32610 9602 32622
rect 9662 32674 9714 32686
rect 9662 32610 9714 32622
rect 16158 32674 16210 32686
rect 22990 32674 23042 32686
rect 18946 32622 18958 32674
rect 19010 32622 19022 32674
rect 20402 32622 20414 32674
rect 20466 32622 20478 32674
rect 16158 32610 16210 32622
rect 22990 32610 23042 32622
rect 23102 32674 23154 32686
rect 23102 32610 23154 32622
rect 25678 32674 25730 32686
rect 25678 32610 25730 32622
rect 30382 32674 30434 32686
rect 30382 32610 30434 32622
rect 30942 32674 30994 32686
rect 30942 32610 30994 32622
rect 32398 32674 32450 32686
rect 32398 32610 32450 32622
rect 32622 32674 32674 32686
rect 32622 32610 32674 32622
rect 34302 32674 34354 32686
rect 34302 32610 34354 32622
rect 39678 32674 39730 32686
rect 39678 32610 39730 32622
rect 39902 32674 39954 32686
rect 39902 32610 39954 32622
rect 40462 32674 40514 32686
rect 40462 32610 40514 32622
rect 5854 32562 5906 32574
rect 14254 32562 14306 32574
rect 1810 32510 1822 32562
rect 1874 32510 1886 32562
rect 13682 32510 13694 32562
rect 13746 32510 13758 32562
rect 5854 32498 5906 32510
rect 14254 32498 14306 32510
rect 14366 32562 14418 32574
rect 15038 32562 15090 32574
rect 14802 32510 14814 32562
rect 14866 32510 14878 32562
rect 14366 32498 14418 32510
rect 15038 32498 15090 32510
rect 15262 32562 15314 32574
rect 15262 32498 15314 32510
rect 15486 32562 15538 32574
rect 15486 32498 15538 32510
rect 15598 32562 15650 32574
rect 15598 32498 15650 32510
rect 16046 32562 16098 32574
rect 16046 32498 16098 32510
rect 16382 32562 16434 32574
rect 18398 32562 18450 32574
rect 17826 32510 17838 32562
rect 17890 32510 17902 32562
rect 16382 32498 16434 32510
rect 18398 32498 18450 32510
rect 18510 32562 18562 32574
rect 21198 32562 21250 32574
rect 18834 32510 18846 32562
rect 18898 32510 18910 32562
rect 19842 32510 19854 32562
rect 19906 32510 19918 32562
rect 18510 32498 18562 32510
rect 21198 32498 21250 32510
rect 23550 32562 23602 32574
rect 23550 32498 23602 32510
rect 30494 32562 30546 32574
rect 30494 32498 30546 32510
rect 30830 32562 30882 32574
rect 30830 32498 30882 32510
rect 32286 32562 32338 32574
rect 32286 32498 32338 32510
rect 33742 32562 33794 32574
rect 38782 32562 38834 32574
rect 34514 32510 34526 32562
rect 34578 32510 34590 32562
rect 34738 32510 34750 32562
rect 34802 32510 34814 32562
rect 35298 32510 35310 32562
rect 35362 32510 35374 32562
rect 33742 32498 33794 32510
rect 38782 32498 38834 32510
rect 39230 32562 39282 32574
rect 39230 32498 39282 32510
rect 40910 32562 40962 32574
rect 40910 32498 40962 32510
rect 42926 32562 42978 32574
rect 42926 32498 42978 32510
rect 43150 32562 43202 32574
rect 43150 32498 43202 32510
rect 43598 32562 43650 32574
rect 51090 32510 51102 32562
rect 51154 32510 51166 32562
rect 43598 32498 43650 32510
rect 5406 32450 5458 32462
rect 2482 32398 2494 32450
rect 2546 32398 2558 32450
rect 4610 32398 4622 32450
rect 4674 32398 4686 32450
rect 5406 32386 5458 32398
rect 7086 32450 7138 32462
rect 7086 32386 7138 32398
rect 13022 32450 13074 32462
rect 13022 32386 13074 32398
rect 16830 32450 16882 32462
rect 16830 32386 16882 32398
rect 21646 32450 21698 32462
rect 21646 32386 21698 32398
rect 24670 32450 24722 32462
rect 24670 32386 24722 32398
rect 25566 32450 25618 32462
rect 25566 32386 25618 32398
rect 29934 32450 29986 32462
rect 29934 32386 29986 32398
rect 31502 32450 31554 32462
rect 31502 32386 31554 32398
rect 31950 32450 32002 32462
rect 38110 32450 38162 32462
rect 34402 32398 34414 32450
rect 34466 32398 34478 32450
rect 35970 32398 35982 32450
rect 36034 32398 36046 32450
rect 31950 32386 32002 32398
rect 38110 32386 38162 32398
rect 39454 32450 39506 32462
rect 39454 32386 39506 32398
rect 42590 32450 42642 32462
rect 42590 32386 42642 32398
rect 53006 32450 53058 32462
rect 53006 32386 53058 32398
rect 25454 32338 25506 32350
rect 25454 32274 25506 32286
rect 30382 32338 30434 32350
rect 30382 32274 30434 32286
rect 1344 32170 53648 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 53648 32170
rect 1344 32084 53648 32118
rect 34638 32002 34690 32014
rect 5618 31950 5630 32002
rect 5682 31950 5694 32002
rect 34638 31938 34690 31950
rect 4846 31890 4898 31902
rect 4846 31826 4898 31838
rect 9998 31890 10050 31902
rect 9998 31826 10050 31838
rect 11118 31890 11170 31902
rect 11118 31826 11170 31838
rect 14590 31890 14642 31902
rect 28366 31890 28418 31902
rect 19618 31838 19630 31890
rect 19682 31838 19694 31890
rect 14590 31826 14642 31838
rect 28366 31826 28418 31838
rect 29262 31890 29314 31902
rect 45602 31838 45614 31890
rect 45666 31838 45678 31890
rect 47730 31838 47742 31890
rect 47794 31838 47806 31890
rect 29262 31826 29314 31838
rect 6190 31778 6242 31790
rect 6190 31714 6242 31726
rect 9102 31778 9154 31790
rect 9102 31714 9154 31726
rect 9326 31778 9378 31790
rect 24558 31778 24610 31790
rect 37102 31778 37154 31790
rect 17826 31726 17838 31778
rect 17890 31726 17902 31778
rect 23426 31726 23438 31778
rect 23490 31726 23502 31778
rect 23986 31726 23998 31778
rect 24050 31726 24062 31778
rect 25442 31726 25454 31778
rect 25506 31726 25518 31778
rect 9326 31714 9378 31726
rect 24558 31714 24610 31726
rect 37102 31714 37154 31726
rect 39230 31778 39282 31790
rect 39230 31714 39282 31726
rect 39678 31778 39730 31790
rect 39678 31714 39730 31726
rect 39902 31778 39954 31790
rect 39902 31714 39954 31726
rect 40686 31778 40738 31790
rect 44158 31778 44210 31790
rect 49982 31778 50034 31790
rect 41122 31726 41134 31778
rect 41186 31726 41198 31778
rect 42802 31726 42814 31778
rect 42866 31726 42878 31778
rect 43474 31726 43486 31778
rect 43538 31726 43550 31778
rect 43810 31726 43822 31778
rect 43874 31726 43886 31778
rect 44930 31726 44942 31778
rect 44994 31726 45006 31778
rect 40686 31714 40738 31726
rect 44158 31714 44210 31726
rect 49982 31714 50034 31726
rect 50430 31778 50482 31790
rect 50430 31714 50482 31726
rect 50542 31778 50594 31790
rect 50542 31714 50594 31726
rect 50990 31778 51042 31790
rect 50990 31714 51042 31726
rect 6078 31666 6130 31678
rect 6078 31602 6130 31614
rect 6302 31666 6354 31678
rect 10558 31666 10610 31678
rect 6738 31614 6750 31666
rect 6802 31614 6814 31666
rect 6302 31602 6354 31614
rect 10558 31602 10610 31614
rect 10670 31666 10722 31678
rect 38894 31666 38946 31678
rect 51214 31666 51266 31678
rect 23650 31614 23662 31666
rect 23714 31614 23726 31666
rect 26226 31614 26238 31666
rect 26290 31614 26302 31666
rect 10670 31602 10722 31614
rect 34638 31610 34690 31622
rect 7086 31554 7138 31566
rect 7086 31490 7138 31502
rect 8878 31554 8930 31566
rect 8878 31490 8930 31502
rect 9214 31554 9266 31566
rect 9214 31490 9266 31502
rect 9774 31554 9826 31566
rect 9774 31490 9826 31502
rect 9886 31554 9938 31566
rect 9886 31490 9938 31502
rect 10334 31554 10386 31566
rect 10334 31490 10386 31502
rect 20302 31554 20354 31566
rect 20302 31490 20354 31502
rect 24222 31554 24274 31566
rect 24222 31490 24274 31502
rect 24334 31554 24386 31566
rect 24334 31490 24386 31502
rect 24446 31554 24498 31566
rect 24446 31490 24498 31502
rect 25118 31554 25170 31566
rect 25118 31490 25170 31502
rect 31950 31554 32002 31566
rect 31950 31490 32002 31502
rect 33742 31554 33794 31566
rect 34638 31546 34690 31558
rect 34750 31610 34802 31622
rect 40226 31614 40238 31666
rect 40290 31614 40302 31666
rect 42690 31614 42702 31666
rect 42754 31614 42766 31666
rect 49074 31614 49086 31666
rect 49138 31614 49150 31666
rect 38894 31602 38946 31614
rect 51214 31602 51266 31614
rect 34750 31546 34802 31558
rect 35198 31554 35250 31566
rect 33742 31490 33794 31502
rect 35198 31490 35250 31502
rect 37550 31554 37602 31566
rect 37550 31490 37602 31502
rect 39006 31554 39058 31566
rect 39006 31490 39058 31502
rect 42366 31554 42418 31566
rect 42366 31490 42418 31502
rect 48750 31554 48802 31566
rect 48750 31490 48802 31502
rect 50654 31554 50706 31566
rect 50654 31490 50706 31502
rect 51102 31554 51154 31566
rect 51102 31490 51154 31502
rect 1344 31386 53648 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 50558 31386
rect 50610 31334 50662 31386
rect 50714 31334 50766 31386
rect 50818 31334 53648 31386
rect 1344 31300 53648 31334
rect 6526 31218 6578 31230
rect 6526 31154 6578 31166
rect 7198 31218 7250 31230
rect 33182 31218 33234 31230
rect 7522 31166 7534 31218
rect 7586 31166 7598 31218
rect 7198 31154 7250 31166
rect 33182 31154 33234 31166
rect 35758 31218 35810 31230
rect 35758 31154 35810 31166
rect 36654 31218 36706 31230
rect 36654 31154 36706 31166
rect 38670 31218 38722 31230
rect 38670 31154 38722 31166
rect 38894 31218 38946 31230
rect 38894 31154 38946 31166
rect 39230 31218 39282 31230
rect 39230 31154 39282 31166
rect 42814 31218 42866 31230
rect 42814 31154 42866 31166
rect 43262 31218 43314 31230
rect 43262 31154 43314 31166
rect 43486 31218 43538 31230
rect 43486 31154 43538 31166
rect 43822 31218 43874 31230
rect 43822 31154 43874 31166
rect 44382 31218 44434 31230
rect 49198 31218 49250 31230
rect 48178 31166 48190 31218
rect 48242 31166 48254 31218
rect 44382 31154 44434 31166
rect 49198 31154 49250 31166
rect 49422 31218 49474 31230
rect 49422 31154 49474 31166
rect 6302 31106 6354 31118
rect 6302 31042 6354 31054
rect 10558 31106 10610 31118
rect 10558 31042 10610 31054
rect 18622 31106 18674 31118
rect 18622 31042 18674 31054
rect 26014 31106 26066 31118
rect 26014 31042 26066 31054
rect 37550 31106 37602 31118
rect 37550 31042 37602 31054
rect 37774 31106 37826 31118
rect 37774 31042 37826 31054
rect 43710 31106 43762 31118
rect 44830 31106 44882 31118
rect 44034 31054 44046 31106
rect 44098 31054 44110 31106
rect 43710 31042 43762 31054
rect 44830 31042 44882 31054
rect 45054 31106 45106 31118
rect 51090 31054 51102 31106
rect 51154 31054 51166 31106
rect 45054 31042 45106 31054
rect 6974 30994 7026 31006
rect 6974 30930 7026 30942
rect 9662 30994 9714 31006
rect 9662 30930 9714 30942
rect 9998 30994 10050 31006
rect 9998 30930 10050 30942
rect 10222 30994 10274 31006
rect 16158 30994 16210 31006
rect 24670 30994 24722 31006
rect 25566 30994 25618 31006
rect 36430 30994 36482 31006
rect 37886 30994 37938 31006
rect 11218 30942 11230 30994
rect 11282 30942 11294 30994
rect 15586 30942 15598 30994
rect 15650 30942 15662 30994
rect 17938 30942 17950 30994
rect 18002 30942 18014 30994
rect 25218 30942 25230 30994
rect 25282 30942 25294 30994
rect 25778 30942 25790 30994
rect 25842 30942 25854 30994
rect 29362 30942 29374 30994
rect 29426 30942 29438 30994
rect 36194 30942 36206 30994
rect 36258 30942 36270 30994
rect 36866 30942 36878 30994
rect 36930 30942 36942 30994
rect 10222 30930 10274 30942
rect 16158 30930 16210 30942
rect 24670 30930 24722 30942
rect 25566 30930 25618 30942
rect 36430 30930 36482 30942
rect 37886 30930 37938 30942
rect 37998 30994 38050 31006
rect 37998 30930 38050 30942
rect 38110 30994 38162 31006
rect 38110 30930 38162 30942
rect 38558 30994 38610 31006
rect 38558 30930 38610 30942
rect 39118 30994 39170 31006
rect 39118 30930 39170 30942
rect 43038 30994 43090 31006
rect 43038 30930 43090 30942
rect 44718 30994 44770 31006
rect 48750 30994 48802 31006
rect 47954 30942 47966 30994
rect 48018 30942 48030 30994
rect 50418 30942 50430 30994
rect 50482 30942 50494 30994
rect 44718 30930 44770 30942
rect 48750 30930 48802 30942
rect 6414 30882 6466 30894
rect 6414 30818 6466 30830
rect 9550 30882 9602 30894
rect 9550 30818 9602 30830
rect 10446 30882 10498 30894
rect 16270 30882 16322 30894
rect 12002 30830 12014 30882
rect 12066 30830 12078 30882
rect 14130 30830 14142 30882
rect 14194 30830 14206 30882
rect 10446 30818 10498 30830
rect 16270 30818 16322 30830
rect 16718 30882 16770 30894
rect 25902 30882 25954 30894
rect 18162 30830 18174 30882
rect 18226 30830 18238 30882
rect 16718 30818 16770 30830
rect 25902 30818 25954 30830
rect 26462 30882 26514 30894
rect 35198 30882 35250 30894
rect 30146 30830 30158 30882
rect 30210 30830 30222 30882
rect 32386 30830 32398 30882
rect 32450 30830 32462 30882
rect 26462 30818 26514 30830
rect 35198 30818 35250 30830
rect 36542 30882 36594 30894
rect 36542 30818 36594 30830
rect 48974 30882 49026 30894
rect 48974 30818 49026 30830
rect 49310 30882 49362 30894
rect 53218 30830 53230 30882
rect 53282 30830 53294 30882
rect 49310 30818 49362 30830
rect 39230 30770 39282 30782
rect 39230 30706 39282 30718
rect 1344 30602 53648 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 53648 30602
rect 1344 30516 53648 30550
rect 9438 30434 9490 30446
rect 9438 30370 9490 30382
rect 9550 30434 9602 30446
rect 9550 30370 9602 30382
rect 9886 30434 9938 30446
rect 9886 30370 9938 30382
rect 30830 30434 30882 30446
rect 30830 30370 30882 30382
rect 50206 30434 50258 30446
rect 50206 30370 50258 30382
rect 9774 30322 9826 30334
rect 25118 30322 25170 30334
rect 11106 30270 11118 30322
rect 11170 30270 11182 30322
rect 16258 30270 16270 30322
rect 16322 30270 16334 30322
rect 23874 30270 23886 30322
rect 23938 30270 23950 30322
rect 9774 30258 9826 30270
rect 25118 30258 25170 30270
rect 36990 30322 37042 30334
rect 50418 30270 50430 30322
rect 50482 30270 50494 30322
rect 36990 30258 37042 30270
rect 13806 30210 13858 30222
rect 20526 30210 20578 30222
rect 12786 30158 12798 30210
rect 12850 30158 12862 30210
rect 16370 30158 16382 30210
rect 16434 30158 16446 30210
rect 13806 30146 13858 30158
rect 20526 30146 20578 30158
rect 20862 30210 20914 30222
rect 20862 30146 20914 30158
rect 21198 30210 21250 30222
rect 21198 30146 21250 30158
rect 21534 30210 21586 30222
rect 21534 30146 21586 30158
rect 21870 30210 21922 30222
rect 26238 30210 26290 30222
rect 23986 30158 23998 30210
rect 24050 30158 24062 30210
rect 25554 30158 25566 30210
rect 25618 30158 25630 30210
rect 21870 30146 21922 30158
rect 26238 30146 26290 30158
rect 29374 30210 29426 30222
rect 29374 30146 29426 30158
rect 30942 30210 30994 30222
rect 30942 30146 30994 30158
rect 34638 30210 34690 30222
rect 35534 30210 35586 30222
rect 35074 30158 35086 30210
rect 35138 30158 35150 30210
rect 34638 30146 34690 30158
rect 35534 30146 35586 30158
rect 38222 30210 38274 30222
rect 42590 30210 42642 30222
rect 41346 30158 41358 30210
rect 41410 30158 41422 30210
rect 50530 30158 50542 30210
rect 50594 30158 50606 30210
rect 38222 30146 38274 30158
rect 42590 30146 42642 30158
rect 20638 30098 20690 30110
rect 13458 30046 13470 30098
rect 13522 30046 13534 30098
rect 20638 30034 20690 30046
rect 23326 30098 23378 30110
rect 23326 30034 23378 30046
rect 29710 30098 29762 30110
rect 29710 30034 29762 30046
rect 29822 30098 29874 30110
rect 29822 30034 29874 30046
rect 30046 30098 30098 30110
rect 30046 30034 30098 30046
rect 30270 30098 30322 30110
rect 30270 30034 30322 30046
rect 30494 30098 30546 30110
rect 30494 30034 30546 30046
rect 31278 30098 31330 30110
rect 31278 30034 31330 30046
rect 31838 30098 31890 30110
rect 35870 30098 35922 30110
rect 35298 30046 35310 30098
rect 35362 30046 35374 30098
rect 31838 30034 31890 30046
rect 35870 30034 35922 30046
rect 52222 30098 52274 30110
rect 52222 30034 52274 30046
rect 53230 30098 53282 30110
rect 53230 30034 53282 30046
rect 4958 29986 5010 29998
rect 4958 29922 5010 29934
rect 16270 29986 16322 29998
rect 16270 29922 16322 29934
rect 21422 29986 21474 29998
rect 21422 29922 21474 29934
rect 23550 29986 23602 29998
rect 23550 29922 23602 29934
rect 23774 29986 23826 29998
rect 23774 29922 23826 29934
rect 24558 29986 24610 29998
rect 24558 29922 24610 29934
rect 30718 29986 30770 29998
rect 30718 29922 30770 29934
rect 31166 29986 31218 29998
rect 33966 29986 34018 29998
rect 35758 29986 35810 29998
rect 33618 29934 33630 29986
rect 33682 29934 33694 29986
rect 34290 29934 34302 29986
rect 34354 29934 34366 29986
rect 31166 29922 31218 29934
rect 33966 29922 34018 29934
rect 35758 29922 35810 29934
rect 36430 29986 36482 29998
rect 36430 29922 36482 29934
rect 37550 29986 37602 29998
rect 37550 29922 37602 29934
rect 41134 29986 41186 29998
rect 41134 29922 41186 29934
rect 42030 29986 42082 29998
rect 42030 29922 42082 29934
rect 52894 29986 52946 29998
rect 52894 29922 52946 29934
rect 1344 29818 53648 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 50558 29818
rect 50610 29766 50662 29818
rect 50714 29766 50766 29818
rect 50818 29766 53648 29818
rect 1344 29732 53648 29766
rect 5406 29650 5458 29662
rect 5406 29586 5458 29598
rect 6190 29650 6242 29662
rect 6190 29586 6242 29598
rect 7086 29650 7138 29662
rect 7086 29586 7138 29598
rect 7310 29650 7362 29662
rect 13022 29650 13074 29662
rect 7970 29598 7982 29650
rect 8034 29598 8046 29650
rect 7310 29586 7362 29598
rect 13022 29586 13074 29598
rect 13470 29650 13522 29662
rect 13470 29586 13522 29598
rect 23214 29650 23266 29662
rect 23214 29586 23266 29598
rect 34302 29650 34354 29662
rect 34302 29586 34354 29598
rect 37886 29650 37938 29662
rect 37886 29586 37938 29598
rect 39006 29650 39058 29662
rect 39006 29586 39058 29598
rect 4958 29538 5010 29550
rect 4958 29474 5010 29486
rect 6078 29538 6130 29550
rect 38222 29538 38274 29550
rect 39566 29538 39618 29550
rect 20402 29486 20414 29538
rect 20466 29486 20478 29538
rect 22866 29486 22878 29538
rect 22930 29486 22942 29538
rect 33954 29486 33966 29538
rect 34018 29486 34030 29538
rect 38434 29486 38446 29538
rect 38498 29486 38510 29538
rect 6078 29474 6130 29486
rect 38222 29474 38274 29486
rect 39566 29474 39618 29486
rect 40238 29538 40290 29550
rect 40238 29474 40290 29486
rect 40350 29538 40402 29550
rect 40350 29474 40402 29486
rect 41246 29538 41298 29550
rect 41246 29474 41298 29486
rect 41806 29538 41858 29550
rect 41806 29474 41858 29486
rect 42142 29538 42194 29550
rect 44930 29486 44942 29538
rect 44994 29486 45006 29538
rect 51090 29486 51102 29538
rect 51154 29486 51166 29538
rect 42142 29474 42194 29486
rect 5182 29426 5234 29438
rect 7422 29426 7474 29438
rect 15374 29426 15426 29438
rect 1810 29374 1822 29426
rect 1874 29374 1886 29426
rect 5618 29374 5630 29426
rect 5682 29374 5694 29426
rect 6850 29374 6862 29426
rect 6914 29374 6926 29426
rect 7970 29374 7982 29426
rect 8034 29374 8046 29426
rect 8194 29374 8206 29426
rect 8258 29374 8270 29426
rect 12338 29374 12350 29426
rect 12402 29374 12414 29426
rect 14802 29374 14814 29426
rect 14866 29374 14878 29426
rect 5182 29362 5234 29374
rect 7422 29362 7474 29374
rect 15374 29362 15426 29374
rect 17502 29426 17554 29438
rect 18846 29426 18898 29438
rect 39454 29426 39506 29438
rect 17714 29374 17726 29426
rect 17778 29374 17790 29426
rect 19618 29374 19630 29426
rect 19682 29374 19694 29426
rect 29138 29374 29150 29426
rect 29202 29374 29214 29426
rect 38994 29374 39006 29426
rect 39058 29374 39070 29426
rect 39890 29374 39902 29426
rect 39954 29423 39966 29426
rect 40114 29423 40126 29426
rect 39954 29377 40126 29423
rect 39954 29374 39966 29377
rect 40114 29374 40126 29377
rect 40178 29374 40190 29426
rect 44258 29374 44270 29426
rect 44322 29374 44334 29426
rect 50418 29374 50430 29426
rect 50482 29374 50494 29426
rect 17502 29362 17554 29374
rect 18846 29362 18898 29374
rect 39454 29362 39506 29374
rect 5294 29314 5346 29326
rect 15486 29314 15538 29326
rect 2482 29262 2494 29314
rect 2546 29262 2558 29314
rect 4610 29262 4622 29314
rect 4674 29262 4686 29314
rect 7858 29262 7870 29314
rect 7922 29262 7934 29314
rect 10098 29262 10110 29314
rect 10162 29262 10174 29314
rect 5294 29250 5346 29262
rect 15486 29250 15538 29262
rect 15934 29314 15986 29326
rect 15934 29250 15986 29262
rect 18398 29314 18450 29326
rect 29710 29314 29762 29326
rect 22530 29262 22542 29314
rect 22594 29262 22606 29314
rect 26114 29262 26126 29314
rect 26178 29262 26190 29314
rect 28354 29262 28366 29314
rect 28418 29262 28430 29314
rect 42578 29262 42590 29314
rect 42642 29262 42654 29314
rect 47058 29262 47070 29314
rect 47122 29262 47134 29314
rect 53218 29262 53230 29314
rect 53282 29262 53294 29314
rect 18398 29250 18450 29262
rect 29710 29250 29762 29262
rect 6302 29202 6354 29214
rect 39342 29202 39394 29214
rect 38770 29150 38782 29202
rect 38834 29150 38846 29202
rect 6302 29138 6354 29150
rect 39342 29138 39394 29150
rect 1344 29034 53648 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 53648 29034
rect 1344 28948 53648 28982
rect 2494 28866 2546 28878
rect 2494 28802 2546 28814
rect 2830 28866 2882 28878
rect 2830 28802 2882 28814
rect 5630 28866 5682 28878
rect 5630 28802 5682 28814
rect 5742 28866 5794 28878
rect 5742 28802 5794 28814
rect 5966 28866 6018 28878
rect 5966 28802 6018 28814
rect 10222 28866 10274 28878
rect 10222 28802 10274 28814
rect 11118 28866 11170 28878
rect 11118 28802 11170 28814
rect 11454 28866 11506 28878
rect 11454 28802 11506 28814
rect 19630 28866 19682 28878
rect 25566 28866 25618 28878
rect 25218 28814 25230 28866
rect 25282 28814 25294 28866
rect 19630 28802 19682 28814
rect 25566 28802 25618 28814
rect 29374 28866 29426 28878
rect 42926 28866 42978 28878
rect 38098 28814 38110 28866
rect 38162 28814 38174 28866
rect 40562 28814 40574 28866
rect 40626 28863 40638 28866
rect 41010 28863 41022 28866
rect 40626 28817 41022 28863
rect 40626 28814 40638 28817
rect 41010 28814 41022 28817
rect 41074 28814 41086 28866
rect 29374 28802 29426 28814
rect 42926 28802 42978 28814
rect 19182 28754 19234 28766
rect 19182 28690 19234 28702
rect 21422 28754 21474 28766
rect 21422 28690 21474 28702
rect 25790 28754 25842 28766
rect 25790 28690 25842 28702
rect 26910 28754 26962 28766
rect 26910 28690 26962 28702
rect 27358 28754 27410 28766
rect 39230 28754 39282 28766
rect 35746 28702 35758 28754
rect 35810 28702 35822 28754
rect 27358 28690 27410 28702
rect 39230 28690 39282 28702
rect 40574 28754 40626 28766
rect 40574 28690 40626 28702
rect 41022 28754 41074 28766
rect 41022 28690 41074 28702
rect 43486 28754 43538 28766
rect 43486 28690 43538 28702
rect 46510 28754 46562 28766
rect 50866 28702 50878 28754
rect 50930 28702 50942 28754
rect 46510 28690 46562 28702
rect 3278 28642 3330 28654
rect 3278 28578 3330 28590
rect 4622 28642 4674 28654
rect 7870 28642 7922 28654
rect 11902 28642 11954 28654
rect 17278 28642 17330 28654
rect 6178 28590 6190 28642
rect 6242 28590 6254 28642
rect 9874 28590 9886 28642
rect 9938 28590 9950 28642
rect 16818 28590 16830 28642
rect 16882 28590 16894 28642
rect 4622 28578 4674 28590
rect 7870 28578 7922 28590
rect 11902 28578 11954 28590
rect 17278 28578 17330 28590
rect 17838 28642 17890 28654
rect 17838 28578 17890 28590
rect 20302 28642 20354 28654
rect 20302 28578 20354 28590
rect 20638 28642 20690 28654
rect 20638 28578 20690 28590
rect 24334 28642 24386 28654
rect 24334 28578 24386 28590
rect 24894 28642 24946 28654
rect 30158 28642 30210 28654
rect 26226 28590 26238 28642
rect 26290 28590 26302 28642
rect 29922 28590 29934 28642
rect 29986 28590 29998 28642
rect 24894 28578 24946 28590
rect 30158 28578 30210 28590
rect 30494 28642 30546 28654
rect 30494 28578 30546 28590
rect 36206 28642 36258 28654
rect 36206 28578 36258 28590
rect 37550 28642 37602 28654
rect 37550 28578 37602 28590
rect 37774 28642 37826 28654
rect 37774 28578 37826 28590
rect 39902 28642 39954 28654
rect 44046 28642 44098 28654
rect 46958 28642 47010 28654
rect 41906 28590 41918 28642
rect 41970 28590 41982 28642
rect 42466 28590 42478 28642
rect 42530 28590 42542 28642
rect 42914 28590 42926 28642
rect 42978 28590 42990 28642
rect 44930 28590 44942 28642
rect 44994 28590 45006 28642
rect 39902 28578 39954 28590
rect 44046 28578 44098 28590
rect 46958 28578 47010 28590
rect 47070 28642 47122 28654
rect 48066 28590 48078 28642
rect 48130 28590 48142 28642
rect 47070 28578 47122 28590
rect 2606 28530 2658 28542
rect 2606 28466 2658 28478
rect 11342 28530 11394 28542
rect 11342 28466 11394 28478
rect 17390 28530 17442 28542
rect 17390 28466 17442 28478
rect 19518 28530 19570 28542
rect 19518 28466 19570 28478
rect 19630 28530 19682 28542
rect 19630 28466 19682 28478
rect 20414 28530 20466 28542
rect 20414 28466 20466 28478
rect 30382 28530 30434 28542
rect 45166 28530 45218 28542
rect 31378 28478 31390 28530
rect 31442 28478 31454 28530
rect 41794 28478 41806 28530
rect 41858 28478 41870 28530
rect 30382 28466 30434 28478
rect 45166 28466 45218 28478
rect 47182 28530 47234 28542
rect 48738 28478 48750 28530
rect 48802 28478 48814 28530
rect 47182 28466 47234 28478
rect 4958 28418 5010 28430
rect 10110 28418 10162 28430
rect 29486 28418 29538 28430
rect 8194 28366 8206 28418
rect 8258 28366 8270 28418
rect 26450 28366 26462 28418
rect 26514 28366 26526 28418
rect 4958 28354 5010 28366
rect 10110 28354 10162 28366
rect 29486 28354 29538 28366
rect 29710 28418 29762 28430
rect 29710 28354 29762 28366
rect 30942 28418 30994 28430
rect 30942 28354 30994 28366
rect 31726 28418 31778 28430
rect 39554 28366 39566 28418
rect 39618 28366 39630 28418
rect 47618 28366 47630 28418
rect 47682 28366 47694 28418
rect 31726 28354 31778 28366
rect 1344 28250 53648 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 50558 28250
rect 50610 28198 50662 28250
rect 50714 28198 50766 28250
rect 50818 28198 53648 28250
rect 1344 28164 53648 28198
rect 7310 28082 7362 28094
rect 7310 28018 7362 28030
rect 10446 28082 10498 28094
rect 10446 28018 10498 28030
rect 11566 28082 11618 28094
rect 21870 28082 21922 28094
rect 25342 28082 25394 28094
rect 18834 28030 18846 28082
rect 18898 28030 18910 28082
rect 22194 28030 22206 28082
rect 22258 28030 22270 28082
rect 23986 28030 23998 28082
rect 24050 28030 24062 28082
rect 24210 28030 24222 28082
rect 24274 28030 24286 28082
rect 11566 28018 11618 28030
rect 21870 28018 21922 28030
rect 25342 28018 25394 28030
rect 26910 28082 26962 28094
rect 26910 28018 26962 28030
rect 34078 28082 34130 28094
rect 36430 28082 36482 28094
rect 34738 28030 34750 28082
rect 34802 28030 34814 28082
rect 35634 28030 35646 28082
rect 35698 28030 35710 28082
rect 34078 28018 34130 28030
rect 36430 28018 36482 28030
rect 36542 28082 36594 28094
rect 36542 28018 36594 28030
rect 41358 28082 41410 28094
rect 44942 28082 44994 28094
rect 43362 28030 43374 28082
rect 43426 28030 43438 28082
rect 41358 28018 41410 28030
rect 44942 28018 44994 28030
rect 48302 28082 48354 28094
rect 48302 28018 48354 28030
rect 48862 28082 48914 28094
rect 48862 28018 48914 28030
rect 48974 28082 49026 28094
rect 48974 28018 49026 28030
rect 5630 27970 5682 27982
rect 5630 27906 5682 27918
rect 5742 27970 5794 27982
rect 5742 27906 5794 27918
rect 10782 27970 10834 27982
rect 19966 27970 20018 27982
rect 52894 27970 52946 27982
rect 10994 27918 11006 27970
rect 11058 27918 11070 27970
rect 12674 27918 12686 27970
rect 12738 27918 12750 27970
rect 17490 27918 17502 27970
rect 17554 27918 17566 27970
rect 22978 27918 22990 27970
rect 23042 27918 23054 27970
rect 31826 27918 31838 27970
rect 31890 27918 31902 27970
rect 34290 27918 34302 27970
rect 34354 27918 34366 27970
rect 38770 27918 38782 27970
rect 38834 27918 38846 27970
rect 10782 27906 10834 27918
rect 19966 27906 20018 27918
rect 39790 27914 39842 27926
rect 40226 27918 40238 27970
rect 40290 27918 40302 27970
rect 5406 27858 5458 27870
rect 5406 27794 5458 27806
rect 7422 27858 7474 27870
rect 7422 27794 7474 27806
rect 8990 27858 9042 27870
rect 8990 27794 9042 27806
rect 9662 27858 9714 27870
rect 9662 27794 9714 27806
rect 10110 27858 10162 27870
rect 10110 27794 10162 27806
rect 10334 27858 10386 27870
rect 16718 27858 16770 27870
rect 22542 27858 22594 27870
rect 36318 27858 36370 27870
rect 37662 27858 37714 27870
rect 52894 27906 52946 27918
rect 11554 27806 11566 27858
rect 11618 27806 11630 27858
rect 11890 27806 11902 27858
rect 11954 27806 11966 27858
rect 16146 27806 16158 27858
rect 16210 27806 16222 27858
rect 17378 27806 17390 27858
rect 17442 27806 17454 27858
rect 19394 27806 19406 27858
rect 19458 27806 19470 27858
rect 23426 27806 23438 27858
rect 23490 27806 23502 27858
rect 23762 27806 23774 27858
rect 23826 27806 23838 27858
rect 27234 27806 27246 27858
rect 27298 27806 27310 27858
rect 34738 27806 34750 27858
rect 34802 27806 34814 27858
rect 35746 27806 35758 27858
rect 35810 27806 35822 27858
rect 36082 27806 36094 27858
rect 36146 27806 36158 27858
rect 36754 27806 36766 27858
rect 36818 27806 36830 27858
rect 38994 27806 39006 27858
rect 39058 27806 39070 27858
rect 39790 27850 39842 27862
rect 53230 27858 53282 27870
rect 40002 27806 40014 27858
rect 40066 27806 40078 27858
rect 10334 27794 10386 27806
rect 16718 27794 16770 27806
rect 22542 27794 22594 27806
rect 36318 27794 36370 27806
rect 37662 27794 37714 27806
rect 53230 27794 53282 27806
rect 8878 27746 8930 27758
rect 16830 27746 16882 27758
rect 14802 27694 14814 27746
rect 14866 27694 14878 27746
rect 8878 27682 8930 27694
rect 16830 27682 16882 27694
rect 26238 27746 26290 27758
rect 26238 27682 26290 27694
rect 37214 27746 37266 27758
rect 37214 27682 37266 27694
rect 43710 27746 43762 27758
rect 43710 27682 43762 27694
rect 43934 27746 43986 27758
rect 43934 27682 43986 27694
rect 44494 27746 44546 27758
rect 44494 27682 44546 27694
rect 45502 27746 45554 27758
rect 45502 27682 45554 27694
rect 52670 27746 52722 27758
rect 52670 27682 52722 27694
rect 9550 27634 9602 27646
rect 9550 27570 9602 27582
rect 11230 27634 11282 27646
rect 48750 27634 48802 27646
rect 44146 27582 44158 27634
rect 44210 27631 44222 27634
rect 44482 27631 44494 27634
rect 44210 27585 44494 27631
rect 44210 27582 44222 27585
rect 44482 27582 44494 27585
rect 44546 27631 44558 27634
rect 44930 27631 44942 27634
rect 44546 27585 44942 27631
rect 44546 27582 44558 27585
rect 44930 27582 44942 27585
rect 44994 27582 45006 27634
rect 11230 27570 11282 27582
rect 48750 27570 48802 27582
rect 1344 27466 53648 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 53648 27466
rect 1344 27380 53648 27414
rect 5966 27298 6018 27310
rect 5966 27234 6018 27246
rect 6190 27298 6242 27310
rect 6190 27234 6242 27246
rect 29262 27298 29314 27310
rect 29262 27234 29314 27246
rect 29822 27298 29874 27310
rect 29822 27234 29874 27246
rect 44270 27298 44322 27310
rect 44270 27234 44322 27246
rect 5070 27186 5122 27198
rect 4610 27134 4622 27186
rect 4674 27134 4686 27186
rect 5070 27122 5122 27134
rect 6414 27186 6466 27198
rect 6414 27122 6466 27134
rect 10670 27186 10722 27198
rect 10670 27122 10722 27134
rect 11790 27186 11842 27198
rect 11790 27122 11842 27134
rect 17166 27186 17218 27198
rect 30606 27186 30658 27198
rect 33966 27186 34018 27198
rect 39790 27186 39842 27198
rect 24658 27134 24670 27186
rect 24722 27134 24734 27186
rect 31826 27134 31838 27186
rect 31890 27134 31902 27186
rect 35298 27134 35310 27186
rect 35362 27134 35374 27186
rect 42018 27134 42030 27186
rect 42082 27134 42094 27186
rect 17166 27122 17218 27134
rect 30606 27122 30658 27134
rect 33966 27122 34018 27134
rect 39790 27122 39842 27134
rect 7086 27074 7138 27086
rect 10446 27074 10498 27086
rect 1810 27022 1822 27074
rect 1874 27022 1886 27074
rect 10210 27022 10222 27074
rect 10274 27022 10286 27074
rect 7086 27010 7138 27022
rect 10446 27010 10498 27022
rect 10782 27074 10834 27086
rect 10782 27010 10834 27022
rect 11118 27074 11170 27086
rect 11118 27010 11170 27022
rect 19070 27074 19122 27086
rect 19070 27010 19122 27022
rect 19630 27074 19682 27086
rect 19630 27010 19682 27022
rect 19966 27074 20018 27086
rect 19966 27010 20018 27022
rect 20190 27074 20242 27086
rect 25006 27074 25058 27086
rect 23314 27022 23326 27074
rect 23378 27022 23390 27074
rect 24210 27022 24222 27074
rect 24274 27022 24286 27074
rect 20190 27010 20242 27022
rect 25006 27010 25058 27022
rect 25342 27074 25394 27086
rect 25342 27010 25394 27022
rect 25790 27074 25842 27086
rect 25790 27010 25842 27022
rect 29374 27074 29426 27086
rect 29374 27010 29426 27022
rect 29934 27074 29986 27086
rect 41470 27074 41522 27086
rect 43934 27074 43986 27086
rect 31154 27022 31166 27074
rect 31218 27022 31230 27074
rect 34626 27022 34638 27074
rect 34690 27022 34702 27074
rect 35746 27022 35758 27074
rect 35810 27022 35822 27074
rect 39330 27022 39342 27074
rect 39394 27022 39406 27074
rect 42130 27022 42142 27074
rect 42194 27022 42206 27074
rect 42466 27022 42478 27074
rect 42530 27022 42542 27074
rect 43698 27022 43710 27074
rect 43762 27022 43774 27074
rect 29934 27010 29986 27022
rect 41470 27010 41522 27022
rect 43934 27010 43986 27022
rect 44158 27074 44210 27086
rect 44158 27010 44210 27022
rect 9774 26962 9826 26974
rect 2482 26910 2494 26962
rect 2546 26910 2558 26962
rect 6738 26910 6750 26962
rect 6802 26910 6814 26962
rect 9774 26898 9826 26910
rect 9998 26962 10050 26974
rect 9998 26898 10050 26910
rect 12238 26962 12290 26974
rect 12238 26898 12290 26910
rect 18958 26962 19010 26974
rect 18958 26898 19010 26910
rect 19294 26962 19346 26974
rect 19294 26898 19346 26910
rect 19406 26962 19458 26974
rect 19406 26898 19458 26910
rect 22990 26962 23042 26974
rect 22990 26898 23042 26910
rect 23550 26962 23602 26974
rect 25230 26962 25282 26974
rect 24322 26910 24334 26962
rect 24386 26910 24398 26962
rect 23550 26898 23602 26910
rect 25230 26898 25282 26910
rect 28590 26962 28642 26974
rect 28590 26898 28642 26910
rect 29262 26962 29314 26974
rect 29262 26898 29314 26910
rect 29822 26962 29874 26974
rect 29822 26898 29874 26910
rect 30270 26962 30322 26974
rect 30270 26898 30322 26910
rect 30718 26962 30770 26974
rect 40238 26962 40290 26974
rect 34738 26910 34750 26962
rect 34802 26910 34814 26962
rect 30718 26898 30770 26910
rect 40238 26898 40290 26910
rect 43374 26962 43426 26974
rect 43374 26898 43426 26910
rect 5518 26850 5570 26862
rect 5518 26786 5570 26798
rect 9662 26850 9714 26862
rect 9662 26786 9714 26798
rect 19854 26850 19906 26862
rect 19854 26786 19906 26798
rect 30494 26850 30546 26862
rect 30494 26786 30546 26798
rect 35870 26850 35922 26862
rect 35870 26786 35922 26798
rect 1344 26682 53648 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 50558 26682
rect 50610 26630 50662 26682
rect 50714 26630 50766 26682
rect 50818 26630 53648 26682
rect 1344 26596 53648 26630
rect 29822 26514 29874 26526
rect 21970 26462 21982 26514
rect 22034 26462 22046 26514
rect 25778 26462 25790 26514
rect 25842 26462 25854 26514
rect 29822 26450 29874 26462
rect 30270 26514 30322 26526
rect 30270 26450 30322 26462
rect 30606 26514 30658 26526
rect 30606 26450 30658 26462
rect 34414 26514 34466 26526
rect 34414 26450 34466 26462
rect 34750 26514 34802 26526
rect 34750 26450 34802 26462
rect 35310 26514 35362 26526
rect 35310 26450 35362 26462
rect 35982 26514 36034 26526
rect 35982 26450 36034 26462
rect 36094 26514 36146 26526
rect 36094 26450 36146 26462
rect 41134 26514 41186 26526
rect 41134 26450 41186 26462
rect 42366 26514 42418 26526
rect 42366 26450 42418 26462
rect 5294 26402 5346 26414
rect 5294 26338 5346 26350
rect 5630 26402 5682 26414
rect 5630 26338 5682 26350
rect 7758 26402 7810 26414
rect 29374 26402 29426 26414
rect 8754 26350 8766 26402
rect 8818 26350 8830 26402
rect 19730 26350 19742 26402
rect 19794 26350 19806 26402
rect 7758 26338 7810 26350
rect 29374 26338 29426 26350
rect 30830 26402 30882 26414
rect 30830 26338 30882 26350
rect 30942 26402 30994 26414
rect 30942 26338 30994 26350
rect 31502 26402 31554 26414
rect 31502 26338 31554 26350
rect 38894 26402 38946 26414
rect 38894 26338 38946 26350
rect 41022 26402 41074 26414
rect 41022 26338 41074 26350
rect 43710 26402 43762 26414
rect 43710 26338 43762 26350
rect 5854 26290 5906 26302
rect 5854 26226 5906 26238
rect 6302 26290 6354 26302
rect 6302 26226 6354 26238
rect 8094 26290 8146 26302
rect 8094 26226 8146 26238
rect 8430 26290 8482 26302
rect 36206 26290 36258 26302
rect 19058 26238 19070 26290
rect 19122 26238 19134 26290
rect 28802 26238 28814 26290
rect 28866 26238 28878 26290
rect 29586 26238 29598 26290
rect 29650 26238 29662 26290
rect 35746 26238 35758 26290
rect 35810 26238 35822 26290
rect 8430 26226 8482 26238
rect 36206 26226 36258 26238
rect 36318 26290 36370 26302
rect 36318 26226 36370 26238
rect 38782 26290 38834 26302
rect 38782 26226 38834 26238
rect 43262 26290 43314 26302
rect 49422 26290 49474 26302
rect 45042 26238 45054 26290
rect 45106 26238 45118 26290
rect 43262 26226 43314 26238
rect 49422 26226 49474 26238
rect 49646 26290 49698 26302
rect 49646 26226 49698 26238
rect 49870 26290 49922 26302
rect 50418 26238 50430 26290
rect 50482 26238 50494 26290
rect 49870 26226 49922 26238
rect 5406 26178 5458 26190
rect 29486 26178 29538 26190
rect 28018 26126 28030 26178
rect 28082 26126 28094 26178
rect 5406 26114 5458 26126
rect 29486 26114 29538 26126
rect 42926 26178 42978 26190
rect 49534 26178 49586 26190
rect 45826 26126 45838 26178
rect 45890 26126 45902 26178
rect 47954 26126 47966 26178
rect 48018 26126 48030 26178
rect 51090 26126 51102 26178
rect 51154 26126 51166 26178
rect 53218 26126 53230 26178
rect 53282 26126 53294 26178
rect 42926 26114 42978 26126
rect 49534 26114 49586 26126
rect 38894 26066 38946 26078
rect 38894 26002 38946 26014
rect 41246 26066 41298 26078
rect 41246 26002 41298 26014
rect 1344 25898 53648 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 53648 25898
rect 1344 25812 53648 25846
rect 29710 25730 29762 25742
rect 45726 25730 45778 25742
rect 31378 25678 31390 25730
rect 31442 25727 31454 25730
rect 31714 25727 31726 25730
rect 31442 25681 31726 25727
rect 31442 25678 31454 25681
rect 31714 25678 31726 25681
rect 31778 25678 31790 25730
rect 29710 25666 29762 25678
rect 45726 25666 45778 25678
rect 50990 25730 51042 25742
rect 50990 25666 51042 25678
rect 29262 25618 29314 25630
rect 17042 25566 17054 25618
rect 17106 25566 17118 25618
rect 24210 25566 24222 25618
rect 24274 25566 24286 25618
rect 26338 25566 26350 25618
rect 26402 25566 26414 25618
rect 29262 25554 29314 25566
rect 31726 25618 31778 25630
rect 37998 25618 38050 25630
rect 37090 25566 37102 25618
rect 37154 25566 37166 25618
rect 31726 25554 31778 25566
rect 37998 25554 38050 25566
rect 42030 25618 42082 25630
rect 45502 25618 45554 25630
rect 42578 25566 42590 25618
rect 42642 25566 42654 25618
rect 42030 25554 42082 25566
rect 45502 25554 45554 25566
rect 49758 25618 49810 25630
rect 49758 25554 49810 25566
rect 51102 25618 51154 25630
rect 51102 25554 51154 25566
rect 7646 25506 7698 25518
rect 7646 25442 7698 25454
rect 7982 25506 8034 25518
rect 10558 25506 10610 25518
rect 8530 25454 8542 25506
rect 8594 25454 8606 25506
rect 9426 25454 9438 25506
rect 9490 25454 9502 25506
rect 7982 25442 8034 25454
rect 10558 25442 10610 25454
rect 10782 25506 10834 25518
rect 10782 25442 10834 25454
rect 11006 25506 11058 25518
rect 11006 25442 11058 25454
rect 11118 25506 11170 25518
rect 11118 25442 11170 25454
rect 11566 25506 11618 25518
rect 19182 25506 19234 25518
rect 16258 25454 16270 25506
rect 16322 25454 16334 25506
rect 11566 25442 11618 25454
rect 19182 25442 19234 25454
rect 19854 25506 19906 25518
rect 19854 25442 19906 25454
rect 23886 25506 23938 25518
rect 30830 25506 30882 25518
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 25554 25454 25566 25506
rect 25618 25454 25630 25506
rect 26226 25454 26238 25506
rect 26290 25454 26302 25506
rect 23886 25442 23938 25454
rect 30830 25442 30882 25454
rect 35422 25506 35474 25518
rect 43150 25506 43202 25518
rect 38994 25454 39006 25506
rect 39058 25454 39070 25506
rect 39778 25454 39790 25506
rect 39842 25454 39854 25506
rect 41122 25454 41134 25506
rect 41186 25454 41198 25506
rect 41570 25454 41582 25506
rect 41634 25454 41646 25506
rect 43026 25454 43038 25506
rect 43090 25454 43102 25506
rect 35422 25442 35474 25454
rect 43150 25442 43202 25454
rect 45838 25506 45890 25518
rect 45838 25442 45890 25454
rect 46062 25506 46114 25518
rect 47742 25506 47794 25518
rect 46274 25454 46286 25506
rect 46338 25454 46350 25506
rect 46062 25442 46114 25454
rect 47742 25442 47794 25454
rect 49870 25506 49922 25518
rect 49870 25442 49922 25454
rect 7198 25394 7250 25406
rect 7198 25330 7250 25342
rect 8094 25394 8146 25406
rect 25230 25394 25282 25406
rect 29822 25394 29874 25406
rect 8194 25342 8206 25394
rect 8258 25342 8270 25394
rect 16594 25342 16606 25394
rect 16658 25342 16670 25394
rect 17602 25342 17614 25394
rect 17666 25342 17678 25394
rect 26002 25342 26014 25394
rect 26066 25342 26078 25394
rect 8094 25330 8146 25342
rect 25230 25330 25282 25342
rect 29822 25330 29874 25342
rect 31166 25394 31218 25406
rect 48190 25394 48242 25406
rect 39330 25342 39342 25394
rect 39394 25342 39406 25394
rect 39666 25342 39678 25394
rect 39730 25342 39742 25394
rect 31166 25330 31218 25342
rect 48190 25330 48242 25342
rect 48414 25394 48466 25406
rect 48414 25330 48466 25342
rect 48750 25394 48802 25406
rect 48750 25330 48802 25342
rect 49086 25394 49138 25406
rect 49086 25330 49138 25342
rect 49310 25394 49362 25406
rect 49310 25330 49362 25342
rect 49646 25394 49698 25406
rect 49646 25330 49698 25342
rect 50206 25394 50258 25406
rect 50206 25330 50258 25342
rect 53230 25394 53282 25406
rect 53230 25330 53282 25342
rect 6414 25282 6466 25294
rect 6066 25230 6078 25282
rect 6130 25230 6142 25282
rect 6414 25218 6466 25230
rect 9886 25282 9938 25294
rect 11902 25282 11954 25294
rect 11106 25230 11118 25282
rect 11170 25230 11182 25282
rect 9886 25218 9938 25230
rect 11902 25218 11954 25230
rect 19518 25282 19570 25294
rect 19518 25218 19570 25230
rect 19742 25282 19794 25294
rect 19742 25218 19794 25230
rect 20302 25282 20354 25294
rect 20302 25218 20354 25230
rect 29710 25282 29762 25294
rect 29710 25218 29762 25230
rect 30382 25282 30434 25294
rect 30382 25218 30434 25230
rect 31054 25282 31106 25294
rect 31054 25218 31106 25230
rect 37550 25282 37602 25294
rect 37550 25218 37602 25230
rect 38558 25282 38610 25294
rect 42254 25282 42306 25294
rect 40002 25230 40014 25282
rect 40066 25230 40078 25282
rect 38558 25218 38610 25230
rect 42254 25218 42306 25230
rect 44046 25282 44098 25294
rect 44046 25218 44098 25230
rect 48078 25282 48130 25294
rect 48078 25218 48130 25230
rect 48862 25282 48914 25294
rect 48862 25218 48914 25230
rect 51214 25282 51266 25294
rect 51214 25218 51266 25230
rect 52894 25282 52946 25294
rect 52894 25218 52946 25230
rect 1344 25114 53648 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 50558 25114
rect 50610 25062 50662 25114
rect 50714 25062 50766 25114
rect 50818 25062 53648 25114
rect 1344 25028 53648 25062
rect 17502 24946 17554 24958
rect 17502 24882 17554 24894
rect 19742 24946 19794 24958
rect 19742 24882 19794 24894
rect 20526 24946 20578 24958
rect 20526 24882 20578 24894
rect 21086 24946 21138 24958
rect 21086 24882 21138 24894
rect 21870 24946 21922 24958
rect 21870 24882 21922 24894
rect 22318 24946 22370 24958
rect 22318 24882 22370 24894
rect 24670 24946 24722 24958
rect 24670 24882 24722 24894
rect 25790 24946 25842 24958
rect 25790 24882 25842 24894
rect 26798 24946 26850 24958
rect 26798 24882 26850 24894
rect 29150 24946 29202 24958
rect 29150 24882 29202 24894
rect 32174 24946 32226 24958
rect 32174 24882 32226 24894
rect 33294 24946 33346 24958
rect 33294 24882 33346 24894
rect 46174 24946 46226 24958
rect 46174 24882 46226 24894
rect 46286 24946 46338 24958
rect 46286 24882 46338 24894
rect 49310 24946 49362 24958
rect 49310 24882 49362 24894
rect 49534 24946 49586 24958
rect 49534 24882 49586 24894
rect 49870 24946 49922 24958
rect 49870 24882 49922 24894
rect 4734 24834 4786 24846
rect 5406 24834 5458 24846
rect 5058 24782 5070 24834
rect 5122 24782 5134 24834
rect 4734 24770 4786 24782
rect 5406 24770 5458 24782
rect 10670 24834 10722 24846
rect 16830 24834 16882 24846
rect 11890 24782 11902 24834
rect 11954 24782 11966 24834
rect 10670 24770 10722 24782
rect 16830 24770 16882 24782
rect 18958 24834 19010 24846
rect 18958 24770 19010 24782
rect 19518 24834 19570 24846
rect 19518 24770 19570 24782
rect 20638 24834 20690 24846
rect 20638 24770 20690 24782
rect 22206 24834 22258 24846
rect 22206 24770 22258 24782
rect 22878 24834 22930 24846
rect 22878 24770 22930 24782
rect 22990 24834 23042 24846
rect 22990 24770 23042 24782
rect 28926 24834 28978 24846
rect 28926 24770 28978 24782
rect 32286 24834 32338 24846
rect 50094 24834 50146 24846
rect 39218 24782 39230 24834
rect 39282 24782 39294 24834
rect 39890 24782 39902 24834
rect 39954 24782 39966 24834
rect 43250 24782 43262 24834
rect 43314 24782 43326 24834
rect 32286 24770 32338 24782
rect 50094 24770 50146 24782
rect 14478 24722 14530 24734
rect 16718 24722 16770 24734
rect 19854 24722 19906 24734
rect 11106 24670 11118 24722
rect 11170 24670 11182 24722
rect 16146 24670 16158 24722
rect 16210 24670 16222 24722
rect 18050 24670 18062 24722
rect 18114 24670 18126 24722
rect 14478 24658 14530 24670
rect 16718 24658 16770 24670
rect 19854 24658 19906 24670
rect 20078 24722 20130 24734
rect 20078 24658 20130 24670
rect 20302 24722 20354 24734
rect 20302 24658 20354 24670
rect 22654 24722 22706 24734
rect 22654 24658 22706 24670
rect 28814 24722 28866 24734
rect 28814 24658 28866 24670
rect 31166 24722 31218 24734
rect 31166 24658 31218 24670
rect 31390 24722 31442 24734
rect 31390 24658 31442 24670
rect 33182 24722 33234 24734
rect 37102 24722 37154 24734
rect 33842 24670 33854 24722
rect 33906 24670 33918 24722
rect 33182 24658 33234 24670
rect 37102 24658 37154 24670
rect 37774 24722 37826 24734
rect 42254 24722 42306 24734
rect 45726 24722 45778 24734
rect 38546 24670 38558 24722
rect 38610 24670 38622 24722
rect 39442 24670 39454 24722
rect 39506 24670 39518 24722
rect 40002 24670 40014 24722
rect 40066 24670 40078 24722
rect 43474 24670 43486 24722
rect 43538 24670 43550 24722
rect 37774 24658 37826 24670
rect 42254 24658 42306 24670
rect 45726 24658 45778 24670
rect 46398 24722 46450 24734
rect 46398 24658 46450 24670
rect 49646 24722 49698 24734
rect 49646 24658 49698 24670
rect 50206 24722 50258 24734
rect 50206 24658 50258 24670
rect 53230 24722 53282 24734
rect 53230 24658 53282 24670
rect 10110 24610 10162 24622
rect 14366 24610 14418 24622
rect 23438 24610 23490 24622
rect 43934 24610 43986 24622
rect 10770 24558 10782 24610
rect 10834 24558 10846 24610
rect 14018 24558 14030 24610
rect 14082 24558 14094 24610
rect 18386 24558 18398 24610
rect 18450 24558 18462 24610
rect 26226 24558 26238 24610
rect 26290 24558 26302 24610
rect 34514 24558 34526 24610
rect 34578 24558 34590 24610
rect 36642 24558 36654 24610
rect 36706 24558 36718 24610
rect 40226 24558 40238 24610
rect 40290 24558 40302 24610
rect 43138 24558 43150 24610
rect 43202 24558 43214 24610
rect 10110 24546 10162 24558
rect 14366 24546 14418 24558
rect 23438 24546 23490 24558
rect 43934 24546 43986 24558
rect 49086 24610 49138 24622
rect 49086 24546 49138 24558
rect 50654 24610 50706 24622
rect 50654 24546 50706 24558
rect 10446 24498 10498 24510
rect 10446 24434 10498 24446
rect 22318 24498 22370 24510
rect 32174 24498 32226 24510
rect 31714 24446 31726 24498
rect 31778 24446 31790 24498
rect 22318 24434 22370 24446
rect 32174 24434 32226 24446
rect 33294 24498 33346 24510
rect 33294 24434 33346 24446
rect 1344 24330 53648 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 53648 24330
rect 1344 24244 53648 24278
rect 34302 24162 34354 24174
rect 34302 24098 34354 24110
rect 45726 24162 45778 24174
rect 45726 24098 45778 24110
rect 5070 24050 5122 24062
rect 7422 24050 7474 24062
rect 26126 24050 26178 24062
rect 4610 23998 4622 24050
rect 4674 23998 4686 24050
rect 6514 23998 6526 24050
rect 6578 23998 6590 24050
rect 8754 23998 8766 24050
rect 8818 23998 8830 24050
rect 17714 23998 17726 24050
rect 17778 23998 17790 24050
rect 19954 23998 19966 24050
rect 20018 23998 20030 24050
rect 24658 23998 24670 24050
rect 24722 23998 24734 24050
rect 5070 23986 5122 23998
rect 7422 23986 7474 23998
rect 26126 23986 26178 23998
rect 28478 24050 28530 24062
rect 28478 23986 28530 23998
rect 40798 24050 40850 24062
rect 40798 23986 40850 23998
rect 47070 24050 47122 24062
rect 47070 23986 47122 23998
rect 5742 23938 5794 23950
rect 1810 23886 1822 23938
rect 1874 23886 1886 23938
rect 5742 23874 5794 23886
rect 7646 23938 7698 23950
rect 7646 23874 7698 23886
rect 8878 23938 8930 23950
rect 8878 23874 8930 23886
rect 15710 23938 15762 23950
rect 31278 23938 31330 23950
rect 20738 23886 20750 23938
rect 20802 23886 20814 23938
rect 21634 23886 21646 23938
rect 21698 23886 21710 23938
rect 25666 23886 25678 23938
rect 25730 23886 25742 23938
rect 15710 23874 15762 23886
rect 31278 23874 31330 23886
rect 31838 23938 31890 23950
rect 37662 23938 37714 23950
rect 34178 23886 34190 23938
rect 34242 23886 34254 23938
rect 31838 23874 31890 23886
rect 37662 23874 37714 23886
rect 39118 23938 39170 23950
rect 39118 23874 39170 23886
rect 41358 23938 41410 23950
rect 46174 23938 46226 23950
rect 43138 23886 43150 23938
rect 43202 23886 43214 23938
rect 41358 23874 41410 23886
rect 46174 23874 46226 23886
rect 5854 23826 5906 23838
rect 2482 23774 2494 23826
rect 2546 23774 2558 23826
rect 5854 23762 5906 23774
rect 6190 23826 6242 23838
rect 6190 23762 6242 23774
rect 6862 23826 6914 23838
rect 6862 23762 6914 23774
rect 8206 23826 8258 23838
rect 8206 23762 8258 23774
rect 8766 23826 8818 23838
rect 8766 23762 8818 23774
rect 9326 23826 9378 23838
rect 27918 23826 27970 23838
rect 15362 23774 15374 23826
rect 15426 23774 15438 23826
rect 22418 23774 22430 23826
rect 22482 23774 22494 23826
rect 9326 23762 9378 23774
rect 27918 23762 27970 23774
rect 28030 23826 28082 23838
rect 28030 23762 28082 23774
rect 33966 23826 34018 23838
rect 33966 23762 34018 23774
rect 34414 23826 34466 23838
rect 34414 23762 34466 23774
rect 34638 23826 34690 23838
rect 34638 23762 34690 23774
rect 34862 23826 34914 23838
rect 34862 23762 34914 23774
rect 34974 23826 35026 23838
rect 34974 23762 35026 23774
rect 37998 23826 38050 23838
rect 37998 23762 38050 23774
rect 38782 23826 38834 23838
rect 38782 23762 38834 23774
rect 38894 23826 38946 23838
rect 38894 23762 38946 23774
rect 42590 23826 42642 23838
rect 42590 23762 42642 23774
rect 43598 23826 43650 23838
rect 43598 23762 43650 23774
rect 44046 23826 44098 23838
rect 44046 23762 44098 23774
rect 45614 23826 45666 23838
rect 45614 23762 45666 23774
rect 5966 23714 6018 23726
rect 5966 23650 6018 23662
rect 6638 23714 6690 23726
rect 6638 23650 6690 23662
rect 7982 23714 8034 23726
rect 7982 23650 8034 23662
rect 8318 23714 8370 23726
rect 8318 23650 8370 23662
rect 9102 23714 9154 23726
rect 9102 23650 9154 23662
rect 25230 23714 25282 23726
rect 25230 23650 25282 23662
rect 26686 23714 26738 23726
rect 26686 23650 26738 23662
rect 27694 23714 27746 23726
rect 32958 23714 33010 23726
rect 30930 23662 30942 23714
rect 30994 23662 31006 23714
rect 32162 23662 32174 23714
rect 32226 23662 32238 23714
rect 27694 23650 27746 23662
rect 32958 23650 33010 23662
rect 37438 23714 37490 23726
rect 37438 23650 37490 23662
rect 37774 23714 37826 23726
rect 37774 23650 37826 23662
rect 43486 23714 43538 23726
rect 43486 23650 43538 23662
rect 45390 23714 45442 23726
rect 45390 23650 45442 23662
rect 45726 23714 45778 23726
rect 45726 23650 45778 23662
rect 46734 23714 46786 23726
rect 46734 23650 46786 23662
rect 47630 23714 47682 23726
rect 47630 23650 47682 23662
rect 1344 23546 53648 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 50558 23546
rect 50610 23494 50662 23546
rect 50714 23494 50766 23546
rect 50818 23494 53648 23546
rect 1344 23460 53648 23494
rect 2606 23378 2658 23390
rect 2606 23314 2658 23326
rect 4734 23378 4786 23390
rect 4734 23314 4786 23326
rect 5406 23378 5458 23390
rect 5406 23314 5458 23326
rect 5630 23378 5682 23390
rect 5630 23314 5682 23326
rect 9774 23378 9826 23390
rect 12350 23378 12402 23390
rect 10546 23326 10558 23378
rect 10610 23326 10622 23378
rect 9774 23314 9826 23326
rect 12350 23314 12402 23326
rect 19294 23378 19346 23390
rect 19294 23314 19346 23326
rect 22542 23378 22594 23390
rect 22542 23314 22594 23326
rect 31166 23378 31218 23390
rect 31838 23378 31890 23390
rect 31490 23326 31502 23378
rect 31554 23326 31566 23378
rect 31166 23314 31218 23326
rect 31838 23314 31890 23326
rect 35198 23378 35250 23390
rect 35198 23314 35250 23326
rect 48862 23378 48914 23390
rect 48862 23314 48914 23326
rect 49086 23378 49138 23390
rect 49086 23314 49138 23326
rect 2830 23266 2882 23278
rect 2830 23202 2882 23214
rect 4510 23266 4562 23278
rect 4510 23202 4562 23214
rect 4958 23266 5010 23278
rect 4958 23202 5010 23214
rect 5854 23266 5906 23278
rect 5854 23202 5906 23214
rect 6190 23266 6242 23278
rect 6190 23202 6242 23214
rect 7646 23266 7698 23278
rect 7646 23202 7698 23214
rect 9550 23266 9602 23278
rect 34750 23266 34802 23278
rect 41694 23266 41746 23278
rect 30818 23214 30830 23266
rect 30882 23214 30894 23266
rect 37650 23214 37662 23266
rect 37714 23214 37726 23266
rect 39330 23214 39342 23266
rect 39394 23214 39406 23266
rect 39554 23214 39566 23266
rect 39618 23214 39630 23266
rect 9550 23202 9602 23214
rect 34750 23202 34802 23214
rect 41694 23202 41746 23214
rect 42030 23266 42082 23278
rect 42030 23202 42082 23214
rect 49758 23266 49810 23278
rect 49758 23202 49810 23214
rect 6302 23154 6354 23166
rect 6302 23090 6354 23102
rect 7198 23154 7250 23166
rect 7198 23090 7250 23102
rect 7870 23154 7922 23166
rect 8654 23154 8706 23166
rect 8418 23102 8430 23154
rect 8482 23102 8494 23154
rect 7870 23090 7922 23102
rect 8654 23090 8706 23102
rect 9998 23154 10050 23166
rect 22318 23154 22370 23166
rect 10210 23102 10222 23154
rect 10274 23102 10286 23154
rect 10770 23102 10782 23154
rect 10834 23102 10846 23154
rect 12674 23102 12686 23154
rect 12738 23102 12750 23154
rect 9998 23090 10050 23102
rect 22318 23090 22370 23102
rect 22654 23154 22706 23166
rect 22654 23090 22706 23102
rect 22990 23154 23042 23166
rect 36654 23154 36706 23166
rect 39230 23154 39282 23166
rect 26450 23102 26462 23154
rect 26514 23102 26526 23154
rect 38098 23102 38110 23154
rect 38162 23102 38174 23154
rect 38434 23102 38446 23154
rect 38498 23102 38510 23154
rect 22990 23090 23042 23102
rect 36654 23090 36706 23102
rect 39230 23090 39282 23102
rect 40014 23154 40066 23166
rect 48750 23154 48802 23166
rect 42802 23102 42814 23154
rect 42866 23102 42878 23154
rect 43026 23102 43038 23154
rect 43090 23102 43102 23154
rect 44146 23102 44158 23154
rect 44210 23102 44222 23154
rect 45714 23102 45726 23154
rect 45778 23102 45790 23154
rect 40014 23090 40066 23102
rect 48750 23090 48802 23102
rect 49310 23154 49362 23166
rect 49310 23090 49362 23102
rect 49870 23154 49922 23166
rect 50418 23102 50430 23154
rect 50482 23102 50494 23154
rect 49870 23090 49922 23102
rect 3278 23042 3330 23054
rect 2482 22990 2494 23042
rect 2546 22990 2558 23042
rect 3278 22978 3330 22990
rect 5742 23042 5794 23054
rect 5742 22978 5794 22990
rect 7422 23042 7474 23054
rect 7422 22978 7474 22990
rect 8990 23042 9042 23054
rect 8990 22978 9042 22990
rect 9886 23042 9938 23054
rect 9886 22978 9938 22990
rect 11342 23042 11394 23054
rect 20974 23042 21026 23054
rect 13458 22990 13470 23042
rect 13522 22990 13534 23042
rect 15586 22990 15598 23042
rect 15650 22990 15662 23042
rect 11342 22978 11394 22990
rect 20974 22978 21026 22990
rect 26126 23042 26178 23054
rect 37214 23042 37266 23054
rect 27234 22990 27246 23042
rect 27298 22990 27310 23042
rect 29362 22990 29374 23042
rect 29426 22990 29438 23042
rect 26126 22978 26178 22990
rect 37214 22978 37266 22990
rect 42142 23042 42194 23054
rect 45278 23042 45330 23054
rect 49534 23042 49586 23054
rect 42690 22990 42702 23042
rect 42754 22990 42766 23042
rect 44482 22990 44494 23042
rect 44546 22990 44558 23042
rect 47954 22990 47966 23042
rect 48018 22990 48030 23042
rect 51090 22990 51102 23042
rect 51154 22990 51166 23042
rect 53218 22990 53230 23042
rect 53282 22990 53294 23042
rect 42142 22978 42194 22990
rect 45278 22978 45330 22990
rect 49534 22978 49586 22990
rect 5070 22930 5122 22942
rect 5070 22866 5122 22878
rect 8878 22930 8930 22942
rect 34738 22878 34750 22930
rect 34802 22927 34814 22930
rect 35186 22927 35198 22930
rect 34802 22881 35198 22927
rect 34802 22878 34814 22881
rect 35186 22878 35198 22881
rect 35250 22878 35262 22930
rect 42578 22878 42590 22930
rect 42642 22878 42654 22930
rect 8878 22866 8930 22878
rect 1344 22762 53648 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 53648 22762
rect 1344 22676 53648 22710
rect 42814 22594 42866 22606
rect 42814 22530 42866 22542
rect 48862 22594 48914 22606
rect 48862 22530 48914 22542
rect 50878 22594 50930 22606
rect 50878 22530 50930 22542
rect 9214 22482 9266 22494
rect 26462 22482 26514 22494
rect 37998 22482 38050 22494
rect 43262 22482 43314 22494
rect 49534 22482 49586 22494
rect 25106 22430 25118 22482
rect 25170 22430 25182 22482
rect 35858 22430 35870 22482
rect 35922 22430 35934 22482
rect 38658 22430 38670 22482
rect 38722 22430 38734 22482
rect 48066 22430 48078 22482
rect 48130 22430 48142 22482
rect 51090 22430 51102 22482
rect 51154 22430 51166 22482
rect 9214 22418 9266 22430
rect 26462 22418 26514 22430
rect 37998 22418 38050 22430
rect 43262 22418 43314 22430
rect 49534 22418 49586 22430
rect 4734 22370 4786 22382
rect 4734 22306 4786 22318
rect 5630 22370 5682 22382
rect 5630 22306 5682 22318
rect 5854 22370 5906 22382
rect 5854 22306 5906 22318
rect 6078 22370 6130 22382
rect 6078 22306 6130 22318
rect 27918 22370 27970 22382
rect 27918 22306 27970 22318
rect 28254 22370 28306 22382
rect 28254 22306 28306 22318
rect 29150 22370 29202 22382
rect 29150 22306 29202 22318
rect 33966 22370 34018 22382
rect 33966 22306 34018 22318
rect 34190 22370 34242 22382
rect 34190 22306 34242 22318
rect 34638 22370 34690 22382
rect 34638 22306 34690 22318
rect 35086 22370 35138 22382
rect 35086 22306 35138 22318
rect 36990 22370 37042 22382
rect 41246 22370 41298 22382
rect 42478 22370 42530 22382
rect 40338 22318 40350 22370
rect 40402 22318 40414 22370
rect 41682 22318 41694 22370
rect 41746 22318 41758 22370
rect 36990 22306 37042 22318
rect 41246 22306 41298 22318
rect 42478 22306 42530 22318
rect 42702 22370 42754 22382
rect 48974 22370 49026 22382
rect 45714 22318 45726 22370
rect 45778 22318 45790 22370
rect 42702 22306 42754 22318
rect 48974 22306 49026 22318
rect 49310 22370 49362 22382
rect 49310 22306 49362 22318
rect 49870 22370 49922 22382
rect 51202 22318 51214 22370
rect 51266 22318 51278 22370
rect 49870 22306 49922 22318
rect 5070 22258 5122 22270
rect 5070 22194 5122 22206
rect 6638 22258 6690 22270
rect 27694 22258 27746 22270
rect 21410 22206 21422 22258
rect 21474 22206 21486 22258
rect 6638 22194 6690 22206
rect 27694 22194 27746 22206
rect 29374 22258 29426 22270
rect 29374 22194 29426 22206
rect 29486 22258 29538 22270
rect 29486 22194 29538 22206
rect 35422 22258 35474 22270
rect 37326 22258 37378 22270
rect 35522 22206 35534 22258
rect 35586 22206 35598 22258
rect 35422 22194 35474 22206
rect 37326 22194 37378 22206
rect 42366 22258 42418 22270
rect 49758 22258 49810 22270
rect 45378 22206 45390 22258
rect 45442 22206 45454 22258
rect 42366 22194 42418 22206
rect 49758 22194 49810 22206
rect 50206 22258 50258 22270
rect 50206 22194 50258 22206
rect 50430 22258 50482 22270
rect 50430 22194 50482 22206
rect 50542 22258 50594 22270
rect 50542 22194 50594 22206
rect 53230 22258 53282 22270
rect 53230 22194 53282 22206
rect 5742 22146 5794 22158
rect 5742 22082 5794 22094
rect 21758 22146 21810 22158
rect 21758 22082 21810 22094
rect 23998 22146 24050 22158
rect 23998 22082 24050 22094
rect 24334 22146 24386 22158
rect 25566 22146 25618 22158
rect 24658 22094 24670 22146
rect 24722 22094 24734 22146
rect 24334 22082 24386 22094
rect 25566 22082 25618 22094
rect 25902 22146 25954 22158
rect 25902 22082 25954 22094
rect 26910 22146 26962 22158
rect 26910 22082 26962 22094
rect 28030 22146 28082 22158
rect 28030 22082 28082 22094
rect 34078 22146 34130 22158
rect 34078 22082 34130 22094
rect 35310 22146 35362 22158
rect 35310 22082 35362 22094
rect 37102 22146 37154 22158
rect 37102 22082 37154 22094
rect 43822 22146 43874 22158
rect 43822 22082 43874 22094
rect 44270 22146 44322 22158
rect 44270 22082 44322 22094
rect 45054 22146 45106 22158
rect 45054 22082 45106 22094
rect 48862 22146 48914 22158
rect 48862 22082 48914 22094
rect 52894 22146 52946 22158
rect 52894 22082 52946 22094
rect 1344 21978 53648 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 50558 21978
rect 50610 21926 50662 21978
rect 50714 21926 50766 21978
rect 50818 21926 53648 21978
rect 1344 21892 53648 21926
rect 5294 21810 5346 21822
rect 5294 21746 5346 21758
rect 5742 21810 5794 21822
rect 5742 21746 5794 21758
rect 8094 21810 8146 21822
rect 8094 21746 8146 21758
rect 8318 21810 8370 21822
rect 8318 21746 8370 21758
rect 9662 21810 9714 21822
rect 14030 21810 14082 21822
rect 13458 21758 13470 21810
rect 13522 21758 13534 21810
rect 9662 21746 9714 21758
rect 14030 21746 14082 21758
rect 21870 21810 21922 21822
rect 21870 21746 21922 21758
rect 22654 21810 22706 21822
rect 22654 21746 22706 21758
rect 34862 21810 34914 21822
rect 34862 21746 34914 21758
rect 38558 21810 38610 21822
rect 38558 21746 38610 21758
rect 41694 21810 41746 21822
rect 46398 21810 46450 21822
rect 43586 21758 43598 21810
rect 43650 21758 43662 21810
rect 41694 21746 41746 21758
rect 46398 21746 46450 21758
rect 49086 21810 49138 21822
rect 49086 21746 49138 21758
rect 49422 21810 49474 21822
rect 49422 21746 49474 21758
rect 49982 21810 50034 21822
rect 49982 21746 50034 21758
rect 53342 21810 53394 21822
rect 53342 21746 53394 21758
rect 23550 21698 23602 21710
rect 2482 21646 2494 21698
rect 2546 21646 2558 21698
rect 23550 21634 23602 21646
rect 23886 21698 23938 21710
rect 23886 21634 23938 21646
rect 33854 21698 33906 21710
rect 47966 21698 48018 21710
rect 35970 21646 35982 21698
rect 36034 21646 36046 21698
rect 40002 21646 40014 21698
rect 40066 21646 40078 21698
rect 44034 21646 44046 21698
rect 44098 21646 44110 21698
rect 33854 21634 33906 21646
rect 47966 21634 48018 21646
rect 48750 21698 48802 21710
rect 48750 21634 48802 21646
rect 48862 21698 48914 21710
rect 48862 21634 48914 21646
rect 49310 21698 49362 21710
rect 49310 21634 49362 21646
rect 7982 21586 8034 21598
rect 20078 21586 20130 21598
rect 1810 21534 1822 21586
rect 1874 21534 1886 21586
rect 10434 21534 10446 21586
rect 10498 21534 10510 21586
rect 19618 21534 19630 21586
rect 19682 21534 19694 21586
rect 7982 21522 8034 21534
rect 20078 21522 20130 21534
rect 20638 21586 20690 21598
rect 20638 21522 20690 21534
rect 21534 21586 21586 21598
rect 21534 21522 21586 21534
rect 23214 21586 23266 21598
rect 23214 21522 23266 21534
rect 33182 21586 33234 21598
rect 33182 21522 33234 21534
rect 33518 21586 33570 21598
rect 41134 21586 41186 21598
rect 45838 21586 45890 21598
rect 35298 21534 35310 21586
rect 35362 21534 35374 21586
rect 40226 21534 40238 21586
rect 40290 21534 40302 21586
rect 40898 21534 40910 21586
rect 40962 21534 40974 21586
rect 43922 21534 43934 21586
rect 43986 21534 43998 21586
rect 33518 21522 33570 21534
rect 41134 21522 41186 21534
rect 45838 21522 45890 21534
rect 47294 21586 47346 21598
rect 47294 21522 47346 21534
rect 47630 21586 47682 21598
rect 47630 21522 47682 21534
rect 49646 21586 49698 21598
rect 49646 21522 49698 21534
rect 8654 21474 8706 21486
rect 4610 21422 4622 21474
rect 4674 21422 4686 21474
rect 8654 21410 8706 21422
rect 9998 21474 10050 21486
rect 15038 21474 15090 21486
rect 11218 21422 11230 21474
rect 11282 21422 11294 21474
rect 9998 21410 10050 21422
rect 15038 21410 15090 21422
rect 15598 21474 15650 21486
rect 15598 21410 15650 21422
rect 19182 21474 19234 21486
rect 19182 21410 19234 21422
rect 22318 21474 22370 21486
rect 22318 21410 22370 21422
rect 33406 21474 33458 21486
rect 42142 21474 42194 21486
rect 38098 21422 38110 21474
rect 38162 21422 38174 21474
rect 39554 21422 39566 21474
rect 39618 21422 39630 21474
rect 33406 21410 33458 21422
rect 42142 21410 42194 21422
rect 44494 21474 44546 21486
rect 44494 21410 44546 21422
rect 44942 21474 44994 21486
rect 44942 21410 44994 21422
rect 45390 21474 45442 21486
rect 45390 21410 45442 21422
rect 46734 21474 46786 21486
rect 46734 21410 46786 21422
rect 50430 21474 50482 21486
rect 50430 21410 50482 21422
rect 10110 21362 10162 21374
rect 10110 21298 10162 21310
rect 41246 21362 41298 21374
rect 44258 21310 44270 21362
rect 44322 21359 44334 21362
rect 44930 21359 44942 21362
rect 44322 21313 44942 21359
rect 44322 21310 44334 21313
rect 44930 21310 44942 21313
rect 44994 21310 45006 21362
rect 41246 21298 41298 21310
rect 1344 21194 53648 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 53648 21194
rect 1344 21108 53648 21142
rect 7534 21026 7586 21038
rect 7534 20962 7586 20974
rect 10446 21026 10498 21038
rect 10446 20962 10498 20974
rect 42814 21026 42866 21038
rect 42814 20962 42866 20974
rect 14590 20914 14642 20926
rect 20414 20914 20466 20926
rect 18498 20862 18510 20914
rect 18562 20862 18574 20914
rect 14590 20850 14642 20862
rect 20414 20850 20466 20862
rect 29822 20914 29874 20926
rect 39230 20914 39282 20926
rect 43486 20914 43538 20926
rect 31714 20862 31726 20914
rect 31778 20862 31790 20914
rect 33842 20862 33854 20914
rect 33906 20862 33918 20914
rect 41010 20862 41022 20914
rect 41074 20862 41086 20914
rect 29822 20850 29874 20862
rect 39230 20850 39282 20862
rect 43486 20850 43538 20862
rect 45390 20914 45442 20926
rect 45390 20850 45442 20862
rect 49982 20914 50034 20926
rect 49982 20850 50034 20862
rect 9998 20802 10050 20814
rect 14142 20802 14194 20814
rect 19966 20802 20018 20814
rect 10210 20750 10222 20802
rect 10274 20750 10286 20802
rect 10546 20750 10558 20802
rect 10610 20750 10622 20802
rect 14802 20750 14814 20802
rect 14866 20750 14878 20802
rect 15586 20750 15598 20802
rect 15650 20750 15662 20802
rect 19058 20750 19070 20802
rect 19122 20750 19134 20802
rect 9998 20738 10050 20750
rect 14142 20738 14194 20750
rect 19966 20738 20018 20750
rect 22206 20802 22258 20814
rect 22206 20738 22258 20750
rect 27022 20802 27074 20814
rect 27022 20738 27074 20750
rect 27694 20802 27746 20814
rect 27694 20738 27746 20750
rect 27918 20802 27970 20814
rect 27918 20738 27970 20750
rect 28254 20802 28306 20814
rect 28254 20738 28306 20750
rect 28478 20802 28530 20814
rect 28478 20738 28530 20750
rect 29374 20802 29426 20814
rect 29374 20738 29426 20750
rect 30270 20802 30322 20814
rect 30270 20738 30322 20750
rect 30606 20802 30658 20814
rect 43038 20802 43090 20814
rect 30930 20750 30942 20802
rect 30994 20750 31006 20802
rect 41570 20750 41582 20802
rect 41634 20750 41646 20802
rect 30606 20738 30658 20750
rect 43038 20738 43090 20750
rect 43262 20802 43314 20814
rect 43262 20738 43314 20750
rect 45950 20802 46002 20814
rect 45950 20738 46002 20750
rect 46510 20802 46562 20814
rect 46510 20738 46562 20750
rect 7870 20690 7922 20702
rect 7870 20626 7922 20638
rect 13806 20690 13858 20702
rect 13806 20626 13858 20638
rect 14478 20690 14530 20702
rect 14478 20626 14530 20638
rect 15262 20690 15314 20702
rect 19630 20690 19682 20702
rect 16370 20638 16382 20690
rect 16434 20638 16446 20690
rect 18834 20638 18846 20690
rect 18898 20638 18910 20690
rect 15262 20626 15314 20638
rect 19630 20626 19682 20638
rect 27246 20690 27298 20702
rect 27246 20626 27298 20638
rect 29038 20690 29090 20702
rect 44942 20690 44994 20702
rect 43810 20638 43822 20690
rect 43874 20638 43886 20690
rect 29038 20626 29090 20638
rect 44942 20626 44994 20638
rect 7646 20578 7698 20590
rect 7646 20514 7698 20526
rect 10782 20578 10834 20590
rect 27358 20578 27410 20590
rect 21858 20526 21870 20578
rect 21922 20526 21934 20578
rect 10782 20514 10834 20526
rect 27358 20514 27410 20526
rect 28366 20578 28418 20590
rect 28366 20514 28418 20526
rect 29262 20578 29314 20590
rect 29262 20514 29314 20526
rect 30494 20578 30546 20590
rect 30494 20514 30546 20526
rect 42366 20578 42418 20590
rect 42366 20514 42418 20526
rect 44158 20578 44210 20590
rect 44158 20514 44210 20526
rect 44830 20578 44882 20590
rect 44830 20514 44882 20526
rect 46958 20578 47010 20590
rect 46958 20514 47010 20526
rect 47406 20578 47458 20590
rect 47406 20514 47458 20526
rect 1344 20410 53648 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 50558 20410
rect 50610 20358 50662 20410
rect 50714 20358 50766 20410
rect 50818 20358 53648 20410
rect 1344 20324 53648 20358
rect 9886 20242 9938 20254
rect 9886 20178 9938 20190
rect 18846 20242 18898 20254
rect 18846 20178 18898 20190
rect 28366 20242 28418 20254
rect 28366 20178 28418 20190
rect 28478 20242 28530 20254
rect 28478 20178 28530 20190
rect 30046 20242 30098 20254
rect 30046 20178 30098 20190
rect 24782 20130 24834 20142
rect 6850 20078 6862 20130
rect 6914 20078 6926 20130
rect 8642 20078 8654 20130
rect 8706 20078 8718 20130
rect 15138 20078 15150 20130
rect 15202 20078 15214 20130
rect 15810 20078 15822 20130
rect 15874 20078 15886 20130
rect 18498 20078 18510 20130
rect 18562 20078 18574 20130
rect 24782 20066 24834 20078
rect 25790 20130 25842 20142
rect 25790 20066 25842 20078
rect 28142 20130 28194 20142
rect 28142 20066 28194 20078
rect 28702 20130 28754 20142
rect 28702 20066 28754 20078
rect 30606 20130 30658 20142
rect 30606 20066 30658 20078
rect 42702 20130 42754 20142
rect 42702 20066 42754 20078
rect 44718 20130 44770 20142
rect 44718 20066 44770 20078
rect 49758 20130 49810 20142
rect 49758 20066 49810 20078
rect 8990 20018 9042 20030
rect 14926 20018 14978 20030
rect 6402 19966 6414 20018
rect 6466 19966 6478 20018
rect 7074 19966 7086 20018
rect 7138 19966 7150 20018
rect 7298 19966 7310 20018
rect 7362 19966 7374 20018
rect 8306 19966 8318 20018
rect 8370 19966 8382 20018
rect 10098 19966 10110 20018
rect 10162 19966 10174 20018
rect 8990 19954 9042 19966
rect 14926 19954 14978 19966
rect 15486 20018 15538 20030
rect 15486 19954 15538 19966
rect 16158 20018 16210 20030
rect 16158 19954 16210 19966
rect 25230 20018 25282 20030
rect 25230 19954 25282 19966
rect 25566 20018 25618 20030
rect 25566 19954 25618 19966
rect 28030 20018 28082 20030
rect 28030 19954 28082 19966
rect 28814 20018 28866 20030
rect 28814 19954 28866 19966
rect 40126 20018 40178 20030
rect 40126 19954 40178 19966
rect 40350 20018 40402 20030
rect 46286 20018 46338 20030
rect 41346 19966 41358 20018
rect 41410 19966 41422 20018
rect 43698 19966 43710 20018
rect 43762 19966 43774 20018
rect 44146 19966 44158 20018
rect 44210 19966 44222 20018
rect 40350 19954 40402 19966
rect 46286 19954 46338 19966
rect 49198 20018 49250 20030
rect 49198 19954 49250 19966
rect 49534 20018 49586 20030
rect 50418 19966 50430 20018
rect 50482 19966 50494 20018
rect 49534 19954 49586 19966
rect 8094 19906 8146 19918
rect 8094 19842 8146 19854
rect 9774 19906 9826 19918
rect 9774 19842 9826 19854
rect 16606 19906 16658 19918
rect 16606 19842 16658 19854
rect 25342 19906 25394 19918
rect 25342 19842 25394 19854
rect 27694 19906 27746 19918
rect 27694 19842 27746 19854
rect 29262 19906 29314 19918
rect 29262 19842 29314 19854
rect 40910 19906 40962 19918
rect 46846 19906 46898 19918
rect 45490 19854 45502 19906
rect 45554 19854 45566 19906
rect 40910 19842 40962 19854
rect 46846 19842 46898 19854
rect 49646 19906 49698 19918
rect 51090 19854 51102 19906
rect 51154 19854 51166 19906
rect 53218 19854 53230 19906
rect 53282 19854 53294 19906
rect 49646 19842 49698 19854
rect 7982 19794 8034 19806
rect 39778 19742 39790 19794
rect 39842 19742 39854 19794
rect 7982 19730 8034 19742
rect 1344 19626 53648 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 53648 19626
rect 1344 19540 53648 19574
rect 4958 19458 5010 19470
rect 11454 19458 11506 19470
rect 7074 19406 7086 19458
rect 7138 19406 7150 19458
rect 4958 19394 5010 19406
rect 11454 19394 11506 19406
rect 38446 19458 38498 19470
rect 38446 19394 38498 19406
rect 51102 19458 51154 19470
rect 51102 19394 51154 19406
rect 8542 19346 8594 19358
rect 8542 19282 8594 19294
rect 11230 19346 11282 19358
rect 11230 19282 11282 19294
rect 12014 19346 12066 19358
rect 12014 19282 12066 19294
rect 15374 19346 15426 19358
rect 31166 19346 31218 19358
rect 41694 19346 41746 19358
rect 18610 19294 18622 19346
rect 18674 19294 18686 19346
rect 23986 19294 23998 19346
rect 24050 19294 24062 19346
rect 26114 19294 26126 19346
rect 26178 19294 26190 19346
rect 30818 19294 30830 19346
rect 30882 19294 30894 19346
rect 39442 19294 39454 19346
rect 39506 19294 39518 19346
rect 15374 19282 15426 19294
rect 31166 19282 31218 19294
rect 41694 19282 41746 19294
rect 45950 19346 46002 19358
rect 45950 19282 46002 19294
rect 5630 19234 5682 19246
rect 5630 19170 5682 19182
rect 5854 19234 5906 19246
rect 7982 19234 8034 19246
rect 7074 19182 7086 19234
rect 7138 19182 7150 19234
rect 5854 19170 5906 19182
rect 7982 19170 8034 19182
rect 8990 19234 9042 19246
rect 31502 19234 31554 19246
rect 10994 19182 11006 19234
rect 11058 19182 11070 19234
rect 15698 19182 15710 19234
rect 15762 19182 15774 19234
rect 23202 19182 23214 19234
rect 23266 19182 23278 19234
rect 30482 19182 30494 19234
rect 30546 19182 30558 19234
rect 8990 19170 9042 19182
rect 31502 19170 31554 19182
rect 32174 19234 32226 19246
rect 32174 19170 32226 19182
rect 32510 19234 32562 19246
rect 34302 19234 34354 19246
rect 33282 19182 33294 19234
rect 33346 19182 33358 19234
rect 32510 19170 32562 19182
rect 34302 19170 34354 19182
rect 34862 19234 34914 19246
rect 46286 19234 46338 19246
rect 49534 19234 49586 19246
rect 39778 19182 39790 19234
rect 39842 19182 39854 19234
rect 47954 19182 47966 19234
rect 48018 19182 48030 19234
rect 34862 19170 34914 19182
rect 46286 19170 46338 19182
rect 49534 19170 49586 19182
rect 49758 19234 49810 19246
rect 49758 19170 49810 19182
rect 49982 19234 50034 19246
rect 49982 19170 50034 19182
rect 53230 19234 53282 19246
rect 53230 19170 53282 19182
rect 5070 19122 5122 19134
rect 5070 19058 5122 19070
rect 6526 19122 6578 19134
rect 11566 19122 11618 19134
rect 22766 19122 22818 19134
rect 6738 19070 6750 19122
rect 6802 19070 6814 19122
rect 7634 19070 7646 19122
rect 7698 19070 7710 19122
rect 10098 19070 10110 19122
rect 10162 19070 10174 19122
rect 16482 19070 16494 19122
rect 16546 19070 16558 19122
rect 6526 19058 6578 19070
rect 11566 19058 11618 19070
rect 22766 19058 22818 19070
rect 22878 19122 22930 19134
rect 22878 19058 22930 19070
rect 31614 19122 31666 19134
rect 31614 19058 31666 19070
rect 31838 19122 31890 19134
rect 31838 19058 31890 19070
rect 32846 19122 32898 19134
rect 32846 19058 32898 19070
rect 34638 19122 34690 19134
rect 34638 19058 34690 19070
rect 35198 19122 35250 19134
rect 38670 19122 38722 19134
rect 35298 19070 35310 19122
rect 35362 19070 35374 19122
rect 35198 19058 35250 19070
rect 38670 19058 38722 19070
rect 39118 19122 39170 19134
rect 48526 19122 48578 19134
rect 46610 19070 46622 19122
rect 46674 19070 46686 19122
rect 39118 19058 39170 19070
rect 48526 19058 48578 19070
rect 48862 19122 48914 19134
rect 48862 19058 48914 19070
rect 49198 19122 49250 19134
rect 49198 19058 49250 19070
rect 50206 19122 50258 19134
rect 50206 19058 50258 19070
rect 50318 19122 50370 19134
rect 50318 19058 50370 19070
rect 50766 19122 50818 19134
rect 50766 19058 50818 19070
rect 50990 19122 51042 19134
rect 50990 19058 51042 19070
rect 52894 19122 52946 19134
rect 52894 19058 52946 19070
rect 4958 19010 5010 19022
rect 6638 19010 6690 19022
rect 6178 18958 6190 19010
rect 6242 18958 6254 19010
rect 4958 18946 5010 18958
rect 6638 18946 6690 18958
rect 10446 19010 10498 19022
rect 10446 18946 10498 18958
rect 22318 19010 22370 19022
rect 22318 18946 22370 18958
rect 22542 19010 22594 19022
rect 22542 18946 22594 18958
rect 32622 19010 32674 19022
rect 32622 18946 32674 18958
rect 32734 19010 32786 19022
rect 32734 18946 32786 18958
rect 33966 19010 34018 19022
rect 33966 18946 34018 18958
rect 34414 19010 34466 19022
rect 34414 18946 34466 18958
rect 34974 19010 35026 19022
rect 34974 18946 35026 18958
rect 35086 19010 35138 19022
rect 35086 18946 35138 18958
rect 38558 19010 38610 19022
rect 38558 18946 38610 18958
rect 42142 19010 42194 19022
rect 49310 19010 49362 19022
rect 48178 18958 48190 19010
rect 48242 18958 48254 19010
rect 42142 18946 42194 18958
rect 49310 18946 49362 18958
rect 1344 18842 53648 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 50558 18842
rect 50610 18790 50662 18842
rect 50714 18790 50766 18842
rect 50818 18790 53648 18842
rect 1344 18756 53648 18790
rect 7646 18674 7698 18686
rect 7646 18610 7698 18622
rect 15150 18674 15202 18686
rect 15150 18610 15202 18622
rect 25118 18674 25170 18686
rect 51102 18674 51154 18686
rect 29250 18622 29262 18674
rect 29314 18622 29326 18674
rect 38322 18622 38334 18674
rect 38386 18622 38398 18674
rect 25118 18610 25170 18622
rect 51102 18610 51154 18622
rect 53342 18674 53394 18686
rect 53342 18610 53394 18622
rect 6414 18562 6466 18574
rect 6414 18498 6466 18510
rect 18510 18562 18562 18574
rect 18510 18498 18562 18510
rect 25342 18562 25394 18574
rect 25342 18498 25394 18510
rect 45502 18562 45554 18574
rect 50094 18562 50146 18574
rect 45826 18510 45838 18562
rect 45890 18510 45902 18562
rect 45502 18498 45554 18510
rect 50094 18498 50146 18510
rect 5966 18450 6018 18462
rect 1810 18398 1822 18450
rect 1874 18398 1886 18450
rect 2482 18398 2494 18450
rect 2546 18398 2558 18450
rect 5506 18398 5518 18450
rect 5570 18398 5582 18450
rect 5966 18386 6018 18398
rect 6302 18450 6354 18462
rect 6302 18386 6354 18398
rect 6638 18450 6690 18462
rect 25454 18450 25506 18462
rect 38894 18450 38946 18462
rect 11890 18398 11902 18450
rect 11954 18398 11966 18450
rect 19842 18398 19854 18450
rect 19906 18398 19918 18450
rect 26226 18398 26238 18450
rect 26290 18398 26302 18450
rect 27010 18398 27022 18450
rect 27074 18398 27086 18450
rect 35410 18398 35422 18450
rect 35474 18398 35486 18450
rect 36082 18398 36094 18450
rect 36146 18398 36158 18450
rect 6638 18386 6690 18398
rect 25454 18386 25506 18398
rect 38894 18386 38946 18398
rect 41806 18450 41858 18462
rect 46734 18450 46786 18462
rect 42242 18398 42254 18450
rect 42306 18398 42318 18450
rect 41806 18386 41858 18398
rect 46734 18386 46786 18398
rect 49870 18450 49922 18462
rect 49870 18386 49922 18398
rect 50542 18450 50594 18462
rect 50542 18386 50594 18398
rect 23214 18338 23266 18350
rect 4610 18286 4622 18338
rect 4674 18286 4686 18338
rect 5058 18286 5070 18338
rect 5122 18286 5134 18338
rect 12562 18286 12574 18338
rect 12626 18286 12638 18338
rect 14690 18286 14702 18338
rect 14754 18286 14766 18338
rect 20626 18286 20638 18338
rect 20690 18286 20702 18338
rect 22754 18286 22766 18338
rect 22818 18286 22830 18338
rect 23214 18274 23266 18286
rect 25902 18338 25954 18350
rect 25902 18274 25954 18286
rect 33182 18338 33234 18350
rect 46174 18338 46226 18350
rect 42914 18286 42926 18338
rect 42978 18286 42990 18338
rect 45042 18286 45054 18338
rect 45106 18286 45118 18338
rect 33182 18274 33234 18286
rect 46174 18274 46226 18286
rect 47182 18338 47234 18350
rect 47182 18274 47234 18286
rect 50318 18338 50370 18350
rect 50318 18274 50370 18286
rect 50878 18338 50930 18350
rect 51090 18286 51102 18338
rect 51154 18286 51166 18338
rect 50878 18274 50930 18286
rect 18398 18226 18450 18238
rect 18398 18162 18450 18174
rect 1344 18058 53648 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 53648 18058
rect 1344 17972 53648 18006
rect 34078 17890 34130 17902
rect 34078 17826 34130 17838
rect 15710 17778 15762 17790
rect 6514 17726 6526 17778
rect 6578 17726 6590 17778
rect 15710 17714 15762 17726
rect 21422 17778 21474 17790
rect 36430 17778 36482 17790
rect 30706 17726 30718 17778
rect 30770 17726 30782 17778
rect 21422 17714 21474 17726
rect 36430 17714 36482 17726
rect 49422 17778 49474 17790
rect 49422 17714 49474 17726
rect 6750 17666 6802 17678
rect 6750 17602 6802 17614
rect 21870 17666 21922 17678
rect 21870 17602 21922 17614
rect 29598 17666 29650 17678
rect 33966 17666 34018 17678
rect 37998 17666 38050 17678
rect 30034 17614 30046 17666
rect 30098 17614 30110 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 29598 17602 29650 17614
rect 33966 17602 34018 17614
rect 37998 17602 38050 17614
rect 38110 17666 38162 17678
rect 43262 17666 43314 17678
rect 39106 17614 39118 17666
rect 39170 17614 39182 17666
rect 40450 17614 40462 17666
rect 40514 17614 40526 17666
rect 42242 17614 42254 17666
rect 42306 17614 42318 17666
rect 38110 17602 38162 17614
rect 43262 17602 43314 17614
rect 48526 17666 48578 17678
rect 48526 17602 48578 17614
rect 49310 17666 49362 17678
rect 49310 17602 49362 17614
rect 49870 17666 49922 17678
rect 49870 17602 49922 17614
rect 6414 17554 6466 17566
rect 6290 17502 6302 17554
rect 6354 17502 6366 17554
rect 6414 17490 6466 17502
rect 6526 17554 6578 17566
rect 15150 17554 15202 17566
rect 7970 17502 7982 17554
rect 8034 17502 8046 17554
rect 6526 17490 6578 17502
rect 15150 17490 15202 17502
rect 21310 17554 21362 17566
rect 21310 17490 21362 17502
rect 21646 17554 21698 17566
rect 21646 17490 21698 17502
rect 23550 17554 23602 17566
rect 23550 17490 23602 17502
rect 23662 17554 23714 17566
rect 23662 17490 23714 17502
rect 33406 17554 33458 17566
rect 47630 17554 47682 17566
rect 38546 17502 38558 17554
rect 38610 17502 38622 17554
rect 42018 17502 42030 17554
rect 42082 17502 42094 17554
rect 33406 17490 33458 17502
rect 47630 17490 47682 17502
rect 48190 17554 48242 17566
rect 48190 17490 48242 17502
rect 48302 17554 48354 17566
rect 48302 17490 48354 17502
rect 49646 17554 49698 17566
rect 49646 17490 49698 17502
rect 4846 17442 4898 17454
rect 4846 17378 4898 17390
rect 7646 17442 7698 17454
rect 7646 17378 7698 17390
rect 15262 17442 15314 17454
rect 15262 17378 15314 17390
rect 23326 17442 23378 17454
rect 33518 17442 33570 17454
rect 32946 17390 32958 17442
rect 33010 17390 33022 17442
rect 23326 17378 23378 17390
rect 33518 17378 33570 17390
rect 36318 17442 36370 17454
rect 36318 17378 36370 17390
rect 40014 17442 40066 17454
rect 47742 17442 47794 17454
rect 42914 17390 42926 17442
rect 42978 17390 42990 17442
rect 40014 17378 40066 17390
rect 47742 17378 47794 17390
rect 47966 17442 48018 17454
rect 47966 17378 48018 17390
rect 48862 17442 48914 17454
rect 48862 17378 48914 17390
rect 1344 17274 53648 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 50558 17274
rect 50610 17222 50662 17274
rect 50714 17222 50766 17274
rect 50818 17222 53648 17274
rect 1344 17188 53648 17222
rect 4622 17106 4674 17118
rect 4622 17042 4674 17054
rect 12910 17106 12962 17118
rect 12910 17042 12962 17054
rect 16606 17106 16658 17118
rect 16606 17042 16658 17054
rect 18174 17106 18226 17118
rect 39006 17106 39058 17118
rect 34514 17054 34526 17106
rect 34578 17054 34590 17106
rect 34738 17054 34750 17106
rect 34802 17054 34814 17106
rect 36306 17054 36318 17106
rect 36370 17054 36382 17106
rect 36530 17054 36542 17106
rect 36594 17054 36606 17106
rect 38098 17054 38110 17106
rect 38162 17054 38174 17106
rect 38322 17054 38334 17106
rect 38386 17054 38398 17106
rect 18174 17042 18226 17054
rect 39006 17042 39058 17054
rect 41246 17106 41298 17118
rect 50094 17106 50146 17118
rect 41906 17054 41918 17106
rect 41970 17054 41982 17106
rect 41246 17042 41298 17054
rect 50094 17042 50146 17054
rect 4734 16994 4786 17006
rect 14478 16994 14530 17006
rect 42702 16994 42754 17006
rect 13010 16942 13022 16994
rect 13074 16942 13086 16994
rect 16034 16942 16046 16994
rect 16098 16942 16110 16994
rect 19282 16942 19294 16994
rect 19346 16942 19358 16994
rect 33730 16942 33742 16994
rect 33794 16942 33806 16994
rect 35410 16942 35422 16994
rect 35474 16942 35486 16994
rect 37090 16942 37102 16994
rect 37154 16942 37166 16994
rect 4734 16930 4786 16942
rect 14478 16930 14530 16942
rect 42702 16930 42754 16942
rect 42814 16994 42866 17006
rect 42814 16930 42866 16942
rect 48862 16994 48914 17006
rect 48862 16930 48914 16942
rect 49758 16994 49810 17006
rect 49758 16930 49810 16942
rect 49870 16994 49922 17006
rect 51090 16942 51102 16994
rect 51154 16942 51166 16994
rect 49870 16930 49922 16942
rect 12798 16882 12850 16894
rect 9650 16830 9662 16882
rect 9714 16830 9726 16882
rect 12798 16818 12850 16830
rect 13246 16882 13298 16894
rect 14590 16882 14642 16894
rect 13458 16830 13470 16882
rect 13522 16830 13534 16882
rect 13246 16818 13298 16830
rect 14590 16818 14642 16830
rect 14814 16882 14866 16894
rect 15822 16882 15874 16894
rect 17390 16882 17442 16894
rect 15250 16830 15262 16882
rect 15314 16830 15326 16882
rect 16594 16830 16606 16882
rect 16658 16830 16670 16882
rect 14814 16818 14866 16830
rect 15822 16818 15874 16830
rect 17390 16818 17442 16830
rect 17726 16882 17778 16894
rect 42030 16882 42082 16894
rect 18162 16830 18174 16882
rect 18226 16830 18238 16882
rect 18610 16830 18622 16882
rect 18674 16830 18686 16882
rect 24098 16830 24110 16882
rect 24162 16830 24174 16882
rect 33394 16830 33406 16882
rect 33458 16830 33470 16882
rect 34290 16830 34302 16882
rect 34354 16830 34366 16882
rect 35298 16830 35310 16882
rect 35362 16830 35374 16882
rect 36418 16830 36430 16882
rect 36482 16830 36494 16882
rect 37538 16830 37550 16882
rect 37602 16830 37614 16882
rect 37874 16830 37886 16882
rect 37938 16830 37950 16882
rect 41570 16830 41582 16882
rect 41634 16830 41646 16882
rect 17726 16818 17778 16830
rect 42030 16818 42082 16830
rect 42366 16882 42418 16894
rect 42366 16818 42418 16830
rect 48750 16882 48802 16894
rect 48750 16818 48802 16830
rect 49086 16882 49138 16894
rect 49086 16818 49138 16830
rect 49422 16882 49474 16894
rect 50306 16830 50318 16882
rect 50370 16830 50382 16882
rect 49422 16818 49474 16830
rect 25342 16770 25394 16782
rect 10322 16718 10334 16770
rect 10386 16718 10398 16770
rect 12450 16718 12462 16770
rect 12514 16718 12526 16770
rect 21410 16718 21422 16770
rect 21474 16718 21486 16770
rect 22306 16718 22318 16770
rect 22370 16718 22382 16770
rect 53218 16718 53230 16770
rect 53282 16718 53294 16770
rect 25342 16706 25394 16718
rect 4510 16658 4562 16670
rect 17838 16658 17890 16670
rect 15026 16606 15038 16658
rect 15090 16606 15102 16658
rect 16370 16606 16382 16658
rect 16434 16606 16446 16658
rect 25106 16606 25118 16658
rect 25170 16655 25182 16658
rect 25330 16655 25342 16658
rect 25170 16609 25342 16655
rect 25170 16606 25182 16609
rect 25330 16606 25342 16609
rect 25394 16606 25406 16658
rect 41794 16606 41806 16658
rect 41858 16606 41870 16658
rect 4510 16594 4562 16606
rect 17838 16594 17890 16606
rect 1344 16490 53648 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 53648 16490
rect 1344 16404 53648 16438
rect 6414 16322 6466 16334
rect 11678 16322 11730 16334
rect 10434 16270 10446 16322
rect 10498 16270 10510 16322
rect 6414 16258 6466 16270
rect 11678 16258 11730 16270
rect 15262 16322 15314 16334
rect 15262 16258 15314 16270
rect 16494 16322 16546 16334
rect 16494 16258 16546 16270
rect 32958 16322 33010 16334
rect 32958 16258 33010 16270
rect 5070 16210 5122 16222
rect 4610 16158 4622 16210
rect 4674 16158 4686 16210
rect 5070 16146 5122 16158
rect 18174 16210 18226 16222
rect 18174 16146 18226 16158
rect 21646 16210 21698 16222
rect 26014 16210 26066 16222
rect 25554 16158 25566 16210
rect 25618 16158 25630 16210
rect 40450 16158 40462 16210
rect 40514 16158 40526 16210
rect 44818 16158 44830 16210
rect 44882 16158 44894 16210
rect 21646 16146 21698 16158
rect 26014 16146 26066 16158
rect 6190 16098 6242 16110
rect 1810 16046 1822 16098
rect 1874 16046 1886 16098
rect 5954 16046 5966 16098
rect 6018 16046 6030 16098
rect 6190 16034 6242 16046
rect 7310 16098 7362 16110
rect 7310 16034 7362 16046
rect 7534 16098 7586 16110
rect 7534 16034 7586 16046
rect 7982 16098 8034 16110
rect 7982 16034 8034 16046
rect 9886 16098 9938 16110
rect 11790 16098 11842 16110
rect 17502 16098 17554 16110
rect 32846 16098 32898 16110
rect 10098 16046 10110 16098
rect 10162 16046 10174 16098
rect 10546 16046 10558 16098
rect 10610 16046 10622 16098
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 16706 16046 16718 16098
rect 16770 16046 16782 16098
rect 17714 16046 17726 16098
rect 17778 16046 17790 16098
rect 22642 16046 22654 16098
rect 22706 16046 22718 16098
rect 9886 16034 9938 16046
rect 11790 16034 11842 16046
rect 17502 16034 17554 16046
rect 32846 16034 32898 16046
rect 37998 16098 38050 16110
rect 37998 16034 38050 16046
rect 38558 16098 38610 16110
rect 38558 16034 38610 16046
rect 38670 16098 38722 16110
rect 42590 16098 42642 16110
rect 48190 16098 48242 16110
rect 40002 16046 40014 16098
rect 40066 16046 40078 16098
rect 40786 16046 40798 16098
rect 40850 16046 40862 16098
rect 47730 16046 47742 16098
rect 47794 16046 47806 16098
rect 38670 16034 38722 16046
rect 42590 16034 42642 16046
rect 48190 16034 48242 16046
rect 48862 16098 48914 16110
rect 48862 16034 48914 16046
rect 49646 16098 49698 16110
rect 49646 16034 49698 16046
rect 50206 16098 50258 16110
rect 53106 16046 53118 16098
rect 53170 16046 53182 16098
rect 50206 16034 50258 16046
rect 6526 15986 6578 15998
rect 2482 15934 2494 15986
rect 2546 15934 2558 15986
rect 6526 15922 6578 15934
rect 15374 15986 15426 15998
rect 15374 15922 15426 15934
rect 15598 15986 15650 15998
rect 15598 15922 15650 15934
rect 16942 15986 16994 15998
rect 16942 15922 16994 15934
rect 17390 15986 17442 15998
rect 34862 15986 34914 15998
rect 42926 15986 42978 15998
rect 48638 15986 48690 15998
rect 23426 15934 23438 15986
rect 23490 15934 23502 15986
rect 38322 15934 38334 15986
rect 38386 15934 38398 15986
rect 39666 15934 39678 15986
rect 39730 15934 39742 15986
rect 40674 15934 40686 15986
rect 40738 15934 40750 15986
rect 46946 15934 46958 15986
rect 47010 15934 47022 15986
rect 17390 15922 17442 15934
rect 34862 15922 34914 15934
rect 42926 15922 42978 15934
rect 48638 15922 48690 15934
rect 49870 15986 49922 15998
rect 49870 15922 49922 15934
rect 52894 15986 52946 15998
rect 52894 15922 52946 15934
rect 7422 15874 7474 15886
rect 12686 15874 12738 15886
rect 37102 15874 37154 15886
rect 10210 15822 10222 15874
rect 10274 15822 10286 15874
rect 16482 15822 16494 15874
rect 16546 15822 16558 15874
rect 7422 15810 7474 15822
rect 12686 15810 12738 15822
rect 37102 15810 37154 15822
rect 37774 15874 37826 15886
rect 37774 15810 37826 15822
rect 42814 15874 42866 15886
rect 42814 15810 42866 15822
rect 48526 15874 48578 15886
rect 48526 15810 48578 15822
rect 50094 15874 50146 15886
rect 50094 15810 50146 15822
rect 1344 15706 53648 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 50558 15706
rect 50610 15654 50662 15706
rect 50714 15654 50766 15706
rect 50818 15654 53648 15706
rect 1344 15620 53648 15654
rect 2270 15538 2322 15550
rect 2270 15474 2322 15486
rect 4622 15538 4674 15550
rect 4622 15474 4674 15486
rect 8542 15538 8594 15550
rect 8542 15474 8594 15486
rect 9662 15538 9714 15550
rect 9662 15474 9714 15486
rect 12126 15538 12178 15550
rect 12126 15474 12178 15486
rect 12798 15538 12850 15550
rect 12798 15474 12850 15486
rect 18510 15538 18562 15550
rect 18510 15474 18562 15486
rect 25342 15538 25394 15550
rect 31390 15538 31442 15550
rect 29810 15486 29822 15538
rect 29874 15486 29886 15538
rect 25342 15474 25394 15486
rect 31390 15474 31442 15486
rect 32398 15538 32450 15550
rect 32398 15474 32450 15486
rect 41022 15538 41074 15550
rect 41022 15474 41074 15486
rect 43262 15538 43314 15550
rect 43262 15474 43314 15486
rect 43486 15538 43538 15550
rect 43486 15474 43538 15486
rect 44494 15538 44546 15550
rect 44494 15474 44546 15486
rect 46398 15538 46450 15550
rect 46398 15474 46450 15486
rect 46734 15538 46786 15550
rect 46734 15474 46786 15486
rect 47966 15538 48018 15550
rect 47966 15474 48018 15486
rect 48638 15538 48690 15550
rect 48638 15474 48690 15486
rect 49870 15538 49922 15550
rect 49870 15474 49922 15486
rect 50430 15538 50482 15550
rect 50430 15474 50482 15486
rect 53342 15538 53394 15550
rect 53342 15474 53394 15486
rect 7086 15426 7138 15438
rect 4946 15374 4958 15426
rect 5010 15374 5022 15426
rect 7086 15362 7138 15374
rect 7198 15426 7250 15438
rect 7198 15362 7250 15374
rect 8206 15426 8258 15438
rect 8206 15362 8258 15374
rect 8766 15426 8818 15438
rect 8766 15362 8818 15374
rect 8878 15426 8930 15438
rect 19742 15426 19794 15438
rect 13122 15374 13134 15426
rect 13186 15374 13198 15426
rect 18610 15374 18622 15426
rect 18674 15374 18686 15426
rect 8878 15362 8930 15374
rect 19742 15362 19794 15374
rect 20750 15426 20802 15438
rect 39790 15426 39842 15438
rect 27570 15374 27582 15426
rect 27634 15374 27646 15426
rect 30930 15374 30942 15426
rect 30994 15374 31006 15426
rect 20750 15362 20802 15374
rect 39790 15362 39842 15374
rect 41470 15426 41522 15438
rect 41470 15362 41522 15374
rect 42366 15426 42418 15438
rect 42366 15362 42418 15374
rect 44606 15426 44658 15438
rect 48862 15426 48914 15438
rect 47058 15374 47070 15426
rect 47122 15374 47134 15426
rect 44606 15362 44658 15374
rect 48862 15362 48914 15374
rect 48974 15426 49026 15438
rect 48974 15362 49026 15374
rect 49534 15426 49586 15438
rect 49534 15362 49586 15374
rect 49646 15426 49698 15438
rect 49646 15362 49698 15374
rect 50094 15426 50146 15438
rect 50094 15362 50146 15374
rect 2606 15314 2658 15326
rect 7982 15314 8034 15326
rect 7522 15262 7534 15314
rect 7586 15262 7598 15314
rect 2606 15250 2658 15262
rect 7982 15250 8034 15262
rect 8094 15314 8146 15326
rect 18398 15314 18450 15326
rect 31614 15314 31666 15326
rect 12338 15262 12350 15314
rect 12402 15262 12414 15314
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 19058 15262 19070 15314
rect 19122 15262 19134 15314
rect 24098 15262 24110 15314
rect 24162 15262 24174 15314
rect 26786 15262 26798 15314
rect 26850 15262 26862 15314
rect 30706 15262 30718 15314
rect 30770 15262 30782 15314
rect 8094 15250 8146 15262
rect 18398 15250 18450 15262
rect 31614 15250 31666 15262
rect 31838 15314 31890 15326
rect 42142 15314 42194 15326
rect 34402 15262 34414 15314
rect 34466 15262 34478 15314
rect 36194 15262 36206 15314
rect 36258 15262 36270 15314
rect 36530 15262 36542 15314
rect 36594 15262 36606 15314
rect 36978 15262 36990 15314
rect 37042 15262 37054 15314
rect 37986 15262 37998 15314
rect 38050 15262 38062 15314
rect 41234 15262 41246 15314
rect 41298 15262 41310 15314
rect 31838 15250 31890 15262
rect 42142 15250 42194 15262
rect 42254 15314 42306 15326
rect 42254 15250 42306 15262
rect 42478 15314 42530 15326
rect 42478 15250 42530 15262
rect 42590 15314 42642 15326
rect 42590 15250 42642 15262
rect 43710 15314 43762 15326
rect 50318 15314 50370 15326
rect 44034 15262 44046 15314
rect 44098 15262 44110 15314
rect 43710 15250 43762 15262
rect 50318 15250 50370 15262
rect 50654 15314 50706 15326
rect 50654 15250 50706 15262
rect 16494 15202 16546 15214
rect 15138 15150 15150 15202
rect 15202 15150 15214 15202
rect 16494 15138 16546 15150
rect 18846 15202 18898 15214
rect 26462 15202 26514 15214
rect 22642 15150 22654 15202
rect 22706 15150 22718 15202
rect 18846 15138 18898 15150
rect 26462 15138 26514 15150
rect 31726 15202 31778 15214
rect 31726 15138 31778 15150
rect 33966 15202 34018 15214
rect 43598 15202 43650 15214
rect 34626 15150 34638 15202
rect 34690 15150 34702 15202
rect 38434 15150 38446 15202
rect 38498 15150 38510 15202
rect 33966 15138 34018 15150
rect 43598 15138 43650 15150
rect 44382 15202 44434 15214
rect 44382 15138 44434 15150
rect 7086 15090 7138 15102
rect 7086 15026 7138 15038
rect 20638 15090 20690 15102
rect 39902 15090 39954 15102
rect 38882 15038 38894 15090
rect 38946 15038 38958 15090
rect 20638 15026 20690 15038
rect 39902 15026 39954 15038
rect 40910 15090 40962 15102
rect 40910 15026 40962 15038
rect 1344 14922 53648 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 53648 14922
rect 1344 14836 53648 14870
rect 19070 14754 19122 14766
rect 19070 14690 19122 14702
rect 31502 14754 31554 14766
rect 31502 14690 31554 14702
rect 33070 14754 33122 14766
rect 33070 14690 33122 14702
rect 35646 14754 35698 14766
rect 35646 14690 35698 14702
rect 23326 14642 23378 14654
rect 15026 14590 15038 14642
rect 15090 14590 15102 14642
rect 23326 14578 23378 14590
rect 34750 14642 34802 14654
rect 52670 14642 52722 14654
rect 41122 14590 41134 14642
rect 41186 14590 41198 14642
rect 34750 14578 34802 14590
rect 52670 14578 52722 14590
rect 6974 14530 7026 14542
rect 11342 14530 11394 14542
rect 7522 14478 7534 14530
rect 7586 14478 7598 14530
rect 10434 14478 10446 14530
rect 10498 14478 10510 14530
rect 6974 14466 7026 14478
rect 11342 14466 11394 14478
rect 12014 14530 12066 14542
rect 16606 14530 16658 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 12014 14466 12066 14478
rect 16606 14466 16658 14478
rect 17278 14530 17330 14542
rect 22878 14530 22930 14542
rect 32174 14530 32226 14542
rect 19058 14478 19070 14530
rect 19122 14478 19134 14530
rect 25330 14478 25342 14530
rect 25394 14478 25406 14530
rect 31938 14478 31950 14530
rect 32002 14478 32014 14530
rect 17278 14466 17330 14478
rect 22878 14466 22930 14478
rect 32174 14466 32226 14478
rect 32510 14530 32562 14542
rect 32510 14466 32562 14478
rect 35870 14530 35922 14542
rect 40686 14530 40738 14542
rect 38658 14478 38670 14530
rect 38722 14478 38734 14530
rect 38882 14478 38894 14530
rect 38946 14478 38958 14530
rect 35870 14466 35922 14478
rect 40686 14466 40738 14478
rect 41022 14530 41074 14542
rect 43374 14530 43426 14542
rect 48526 14530 48578 14542
rect 41234 14478 41246 14530
rect 41298 14478 41310 14530
rect 46386 14478 46398 14530
rect 46450 14478 46462 14530
rect 41022 14466 41074 14478
rect 43374 14466 43426 14478
rect 48526 14466 48578 14478
rect 48862 14530 48914 14542
rect 48862 14466 48914 14478
rect 49086 14530 49138 14542
rect 49086 14466 49138 14478
rect 11006 14418 11058 14430
rect 11006 14354 11058 14366
rect 18734 14418 18786 14430
rect 18734 14354 18786 14366
rect 23102 14418 23154 14430
rect 23102 14354 23154 14366
rect 23438 14418 23490 14430
rect 31278 14418 31330 14430
rect 25778 14366 25790 14418
rect 25842 14366 25854 14418
rect 23438 14354 23490 14366
rect 31278 14354 31330 14366
rect 32286 14418 32338 14430
rect 32286 14354 32338 14366
rect 33182 14418 33234 14430
rect 39118 14418 39170 14430
rect 46062 14418 46114 14430
rect 35298 14366 35310 14418
rect 35362 14366 35374 14418
rect 41906 14366 41918 14418
rect 41970 14366 41982 14418
rect 43026 14366 43038 14418
rect 43090 14366 43102 14418
rect 33182 14354 33234 14366
rect 39118 14354 39170 14366
rect 46062 14354 46114 14366
rect 7086 14306 7138 14318
rect 7086 14242 7138 14254
rect 7198 14306 7250 14318
rect 7198 14242 7250 14254
rect 8542 14306 8594 14318
rect 11678 14306 11730 14318
rect 10210 14254 10222 14306
rect 10274 14254 10286 14306
rect 8542 14242 8594 14254
rect 11678 14242 11730 14254
rect 16942 14306 16994 14318
rect 16942 14242 16994 14254
rect 17614 14306 17666 14318
rect 26126 14306 26178 14318
rect 25106 14254 25118 14306
rect 25170 14254 25182 14306
rect 17614 14242 17666 14254
rect 26126 14242 26178 14254
rect 26574 14306 26626 14318
rect 26574 14242 26626 14254
rect 31390 14306 31442 14318
rect 31390 14242 31442 14254
rect 32398 14306 32450 14318
rect 32398 14242 32450 14254
rect 33070 14306 33122 14318
rect 33070 14242 33122 14254
rect 40798 14306 40850 14318
rect 40798 14242 40850 14254
rect 42254 14306 42306 14318
rect 42254 14242 42306 14254
rect 46174 14306 46226 14318
rect 46174 14242 46226 14254
rect 46846 14306 46898 14318
rect 46846 14242 46898 14254
rect 48862 14306 48914 14318
rect 48862 14242 48914 14254
rect 52222 14306 52274 14318
rect 52222 14242 52274 14254
rect 53230 14306 53282 14318
rect 53230 14242 53282 14254
rect 1344 14138 53648 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 50558 14138
rect 50610 14086 50662 14138
rect 50714 14086 50766 14138
rect 50818 14086 53648 14138
rect 1344 14052 53648 14086
rect 7310 13970 7362 13982
rect 10334 13970 10386 13982
rect 15598 13970 15650 13982
rect 9538 13918 9550 13970
rect 9602 13918 9614 13970
rect 12562 13918 12574 13970
rect 12626 13918 12638 13970
rect 7310 13906 7362 13918
rect 10334 13906 10386 13918
rect 15598 13906 15650 13918
rect 16942 13970 16994 13982
rect 32286 13970 32338 13982
rect 18610 13918 18622 13970
rect 18674 13918 18686 13970
rect 16942 13906 16994 13918
rect 32286 13906 32338 13918
rect 33854 13970 33906 13982
rect 33854 13906 33906 13918
rect 39678 13970 39730 13982
rect 40002 13918 40014 13970
rect 40066 13918 40078 13970
rect 39678 13906 39730 13918
rect 16382 13858 16434 13870
rect 16146 13806 16158 13858
rect 16210 13806 16222 13858
rect 16382 13794 16434 13806
rect 18286 13858 18338 13870
rect 18286 13794 18338 13806
rect 19630 13858 19682 13870
rect 31838 13858 31890 13870
rect 27906 13806 27918 13858
rect 27970 13806 27982 13858
rect 19630 13794 19682 13806
rect 31838 13794 31890 13806
rect 32510 13858 32562 13870
rect 32510 13794 32562 13806
rect 33630 13858 33682 13870
rect 33630 13794 33682 13806
rect 5966 13746 6018 13758
rect 5170 13694 5182 13746
rect 5234 13694 5246 13746
rect 5966 13682 6018 13694
rect 6190 13746 6242 13758
rect 6190 13682 6242 13694
rect 6414 13746 6466 13758
rect 6974 13746 7026 13758
rect 15934 13746 15986 13758
rect 20302 13746 20354 13758
rect 32062 13746 32114 13758
rect 6626 13694 6638 13746
rect 6690 13694 6702 13746
rect 9762 13694 9774 13746
rect 9826 13694 9838 13746
rect 12338 13694 12350 13746
rect 12402 13694 12414 13746
rect 15810 13694 15822 13746
rect 15874 13694 15886 13746
rect 18498 13694 18510 13746
rect 18562 13694 18574 13746
rect 19058 13694 19070 13746
rect 19122 13694 19134 13746
rect 21522 13694 21534 13746
rect 21586 13694 21598 13746
rect 27122 13694 27134 13746
rect 27186 13694 27198 13746
rect 35522 13694 35534 13746
rect 35586 13694 35598 13746
rect 50306 13694 50318 13746
rect 50370 13694 50382 13746
rect 6414 13682 6466 13694
rect 6974 13682 7026 13694
rect 15934 13682 15986 13694
rect 20302 13682 20354 13694
rect 32062 13682 32114 13694
rect 6078 13634 6130 13646
rect 5058 13582 5070 13634
rect 5122 13582 5134 13634
rect 6078 13570 6130 13582
rect 17614 13634 17666 13646
rect 17614 13570 17666 13582
rect 18734 13634 18786 13646
rect 18734 13570 18786 13582
rect 19518 13634 19570 13646
rect 25342 13634 25394 13646
rect 22194 13582 22206 13634
rect 22258 13582 22270 13634
rect 24322 13582 24334 13634
rect 24386 13582 24398 13634
rect 19518 13570 19570 13582
rect 25342 13570 25394 13582
rect 26798 13634 26850 13646
rect 36206 13634 36258 13646
rect 30034 13582 30046 13634
rect 30098 13582 30110 13634
rect 35746 13582 35758 13634
rect 35810 13582 35822 13634
rect 26798 13570 26850 13582
rect 36206 13570 36258 13582
rect 49982 13634 50034 13646
rect 51090 13582 51102 13634
rect 51154 13582 51166 13634
rect 53218 13582 53230 13634
rect 53282 13582 53294 13634
rect 49982 13570 50034 13582
rect 4846 13522 4898 13534
rect 19406 13522 19458 13534
rect 7074 13470 7086 13522
rect 7138 13519 7150 13522
rect 7410 13519 7422 13522
rect 7138 13473 7422 13519
rect 7138 13470 7150 13473
rect 7410 13470 7422 13473
rect 7474 13470 7486 13522
rect 4846 13458 4898 13470
rect 19406 13458 19458 13470
rect 31950 13522 32002 13534
rect 31950 13458 32002 13470
rect 33966 13522 34018 13534
rect 33966 13458 34018 13470
rect 1344 13354 53648 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 53648 13354
rect 1344 13268 53648 13302
rect 6190 13186 6242 13198
rect 6190 13122 6242 13134
rect 6414 13186 6466 13198
rect 6414 13122 6466 13134
rect 6862 13186 6914 13198
rect 6862 13122 6914 13134
rect 10670 13186 10722 13198
rect 10670 13122 10722 13134
rect 14366 13186 14418 13198
rect 14366 13122 14418 13134
rect 15486 13186 15538 13198
rect 15486 13122 15538 13134
rect 15822 13186 15874 13198
rect 41918 13186 41970 13198
rect 18610 13134 18622 13186
rect 18674 13134 18686 13186
rect 15822 13122 15874 13134
rect 41918 13122 41970 13134
rect 50542 13186 50594 13198
rect 50542 13122 50594 13134
rect 50878 13186 50930 13198
rect 50878 13122 50930 13134
rect 4958 13074 5010 13086
rect 2482 13022 2494 13074
rect 2546 13022 2558 13074
rect 4610 13022 4622 13074
rect 4674 13022 4686 13074
rect 4958 13010 5010 13022
rect 7198 13074 7250 13086
rect 7198 13010 7250 13022
rect 11566 13074 11618 13086
rect 11566 13010 11618 13022
rect 11902 13074 11954 13086
rect 11902 13010 11954 13022
rect 22206 13074 22258 13086
rect 22206 13010 22258 13022
rect 24782 13074 24834 13086
rect 28578 13022 28590 13074
rect 28642 13022 28654 13074
rect 46834 13022 46846 13074
rect 46898 13022 46910 13074
rect 24782 13010 24834 13022
rect 5070 12962 5122 12974
rect 1810 12910 1822 12962
rect 1874 12910 1886 12962
rect 5070 12898 5122 12910
rect 5742 12962 5794 12974
rect 13918 12962 13970 12974
rect 6850 12910 6862 12962
rect 6914 12910 6926 12962
rect 10994 12910 11006 12962
rect 11058 12910 11070 12962
rect 5742 12898 5794 12910
rect 13918 12898 13970 12910
rect 14254 12962 14306 12974
rect 15150 12962 15202 12974
rect 18062 12962 18114 12974
rect 14466 12910 14478 12962
rect 14530 12910 14542 12962
rect 15810 12910 15822 12962
rect 15874 12910 15886 12962
rect 14254 12898 14306 12910
rect 15150 12898 15202 12910
rect 18062 12898 18114 12910
rect 18398 12962 18450 12974
rect 21870 12962 21922 12974
rect 18834 12910 18846 12962
rect 18898 12910 18910 12962
rect 18398 12898 18450 12910
rect 21870 12898 21922 12910
rect 22094 12962 22146 12974
rect 22094 12898 22146 12910
rect 22430 12962 22482 12974
rect 36206 12962 36258 12974
rect 38334 12962 38386 12974
rect 25666 12910 25678 12962
rect 25730 12910 25742 12962
rect 35634 12910 35646 12962
rect 35698 12910 35710 12962
rect 38098 12910 38110 12962
rect 38162 12910 38174 12962
rect 38770 12910 38782 12962
rect 38834 12910 38846 12962
rect 42242 12910 42254 12962
rect 42306 12910 42318 12962
rect 43922 12910 43934 12962
rect 43986 12910 43998 12962
rect 49746 12910 49758 12962
rect 49810 12910 49822 12962
rect 22430 12898 22482 12910
rect 36206 12898 36258 12910
rect 38334 12898 38386 12910
rect 5630 12850 5682 12862
rect 5630 12786 5682 12798
rect 23998 12850 24050 12862
rect 23998 12786 24050 12798
rect 24222 12850 24274 12862
rect 24222 12786 24274 12798
rect 24334 12850 24386 12862
rect 26450 12798 26462 12850
rect 26514 12798 26526 12850
rect 43698 12798 43710 12850
rect 43762 12798 43774 12850
rect 48962 12798 48974 12850
rect 49026 12798 49038 12850
rect 24334 12786 24386 12798
rect 6526 12738 6578 12750
rect 6526 12674 6578 12686
rect 10782 12738 10834 12750
rect 10782 12674 10834 12686
rect 14702 12738 14754 12750
rect 14702 12674 14754 12686
rect 18174 12738 18226 12750
rect 18174 12674 18226 12686
rect 25342 12738 25394 12750
rect 25342 12674 25394 12686
rect 35870 12738 35922 12750
rect 35870 12674 35922 12686
rect 35982 12738 36034 12750
rect 35982 12674 36034 12686
rect 36094 12738 36146 12750
rect 36094 12674 36146 12686
rect 38446 12738 38498 12750
rect 38446 12674 38498 12686
rect 38558 12738 38610 12750
rect 38558 12674 38610 12686
rect 42030 12738 42082 12750
rect 42030 12674 42082 12686
rect 45614 12738 45666 12750
rect 46286 12738 46338 12750
rect 45938 12686 45950 12738
rect 46002 12686 46014 12738
rect 45614 12674 45666 12686
rect 46286 12674 46338 12686
rect 50206 12738 50258 12750
rect 50206 12674 50258 12686
rect 50766 12738 50818 12750
rect 50766 12674 50818 12686
rect 1344 12570 53648 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 50558 12570
rect 50610 12518 50662 12570
rect 50714 12518 50766 12570
rect 50818 12518 53648 12570
rect 1344 12484 53648 12518
rect 10670 12402 10722 12414
rect 10670 12338 10722 12350
rect 14030 12402 14082 12414
rect 14030 12338 14082 12350
rect 24110 12402 24162 12414
rect 24110 12338 24162 12350
rect 27022 12402 27074 12414
rect 27022 12338 27074 12350
rect 27694 12402 27746 12414
rect 27694 12338 27746 12350
rect 28814 12402 28866 12414
rect 28814 12338 28866 12350
rect 41022 12402 41074 12414
rect 41022 12338 41074 12350
rect 45390 12402 45442 12414
rect 45390 12338 45442 12350
rect 45726 12402 45778 12414
rect 45726 12338 45778 12350
rect 48862 12402 48914 12414
rect 48862 12338 48914 12350
rect 9886 12290 9938 12302
rect 9886 12226 9938 12238
rect 12126 12290 12178 12302
rect 12126 12226 12178 12238
rect 13918 12290 13970 12302
rect 13918 12226 13970 12238
rect 14142 12290 14194 12302
rect 14142 12226 14194 12238
rect 14590 12290 14642 12302
rect 14590 12226 14642 12238
rect 14814 12290 14866 12302
rect 14814 12226 14866 12238
rect 27582 12290 27634 12302
rect 27582 12226 27634 12238
rect 36318 12290 36370 12302
rect 36318 12226 36370 12238
rect 36542 12290 36594 12302
rect 36542 12226 36594 12238
rect 48750 12290 48802 12302
rect 48750 12226 48802 12238
rect 48974 12290 49026 12302
rect 52434 12238 52446 12290
rect 52498 12238 52510 12290
rect 48974 12226 49026 12238
rect 8094 12178 8146 12190
rect 12462 12178 12514 12190
rect 13470 12178 13522 12190
rect 10098 12126 10110 12178
rect 10162 12126 10174 12178
rect 10658 12126 10670 12178
rect 10722 12126 10734 12178
rect 12898 12126 12910 12178
rect 12962 12126 12974 12178
rect 8094 12114 8146 12126
rect 12462 12114 12514 12126
rect 13470 12114 13522 12126
rect 21758 12178 21810 12190
rect 21758 12114 21810 12126
rect 21870 12178 21922 12190
rect 21870 12114 21922 12126
rect 22318 12178 22370 12190
rect 22318 12114 22370 12126
rect 23886 12178 23938 12190
rect 23886 12114 23938 12126
rect 24222 12178 24274 12190
rect 24222 12114 24274 12126
rect 26686 12178 26738 12190
rect 26686 12114 26738 12126
rect 26910 12178 26962 12190
rect 26910 12114 26962 12126
rect 27358 12178 27410 12190
rect 29250 12126 29262 12178
rect 29314 12126 29326 12178
rect 35970 12126 35982 12178
rect 36034 12126 36046 12178
rect 37090 12126 37102 12178
rect 37154 12126 37166 12178
rect 41570 12126 41582 12178
rect 41634 12126 41646 12178
rect 27358 12114 27410 12126
rect 4846 12066 4898 12078
rect 4846 12002 4898 12014
rect 7870 12066 7922 12078
rect 7870 12002 7922 12014
rect 12238 12066 12290 12078
rect 19294 12066 19346 12078
rect 14466 12014 14478 12066
rect 14530 12014 14542 12066
rect 12238 12002 12290 12014
rect 19294 12002 19346 12014
rect 22094 12066 22146 12078
rect 22094 12002 22146 12014
rect 24670 12066 24722 12078
rect 36430 12066 36482 12078
rect 52782 12066 52834 12078
rect 29922 12014 29934 12066
rect 29986 12014 29998 12066
rect 32050 12014 32062 12066
rect 32114 12014 32126 12066
rect 33058 12014 33070 12066
rect 33122 12014 33134 12066
rect 35186 12014 35198 12066
rect 35250 12014 35262 12066
rect 37874 12014 37886 12066
rect 37938 12014 37950 12066
rect 40002 12014 40014 12066
rect 40066 12014 40078 12066
rect 42354 12014 42366 12066
rect 42418 12014 42430 12066
rect 44482 12014 44494 12066
rect 44546 12014 44558 12066
rect 46162 12014 46174 12066
rect 46226 12014 46238 12066
rect 24670 12002 24722 12014
rect 36430 12002 36482 12014
rect 52782 12002 52834 12014
rect 53342 12066 53394 12078
rect 53342 12002 53394 12014
rect 8318 11954 8370 11966
rect 8318 11890 8370 11902
rect 8766 11954 8818 11966
rect 8766 11890 8818 11902
rect 10334 11954 10386 11966
rect 10334 11890 10386 11902
rect 12574 11954 12626 11966
rect 12574 11890 12626 11902
rect 19182 11954 19234 11966
rect 19182 11890 19234 11902
rect 27694 11954 27746 11966
rect 27694 11890 27746 11902
rect 1344 11786 53648 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 53648 11786
rect 1344 11700 53648 11734
rect 15598 11618 15650 11630
rect 15598 11554 15650 11566
rect 38110 11618 38162 11630
rect 38110 11554 38162 11566
rect 38446 11618 38498 11630
rect 40450 11566 40462 11618
rect 40514 11615 40526 11618
rect 41010 11615 41022 11618
rect 40514 11569 41022 11615
rect 40514 11566 40526 11569
rect 41010 11566 41022 11569
rect 41074 11566 41086 11618
rect 42018 11566 42030 11618
rect 42082 11566 42094 11618
rect 38446 11554 38498 11566
rect 5854 11506 5906 11518
rect 5854 11442 5906 11454
rect 7870 11506 7922 11518
rect 7870 11442 7922 11454
rect 14478 11506 14530 11518
rect 31838 11506 31890 11518
rect 17714 11454 17726 11506
rect 17778 11454 17790 11506
rect 19842 11454 19854 11506
rect 19906 11454 19918 11506
rect 22194 11454 22206 11506
rect 22258 11454 22270 11506
rect 24322 11454 24334 11506
rect 24386 11454 24398 11506
rect 14478 11442 14530 11454
rect 31838 11442 31890 11454
rect 41246 11506 41298 11518
rect 41246 11442 41298 11454
rect 42478 11506 42530 11518
rect 42478 11442 42530 11454
rect 6078 11394 6130 11406
rect 6638 11394 6690 11406
rect 6290 11342 6302 11394
rect 6354 11342 6366 11394
rect 6078 11330 6130 11342
rect 6638 11330 6690 11342
rect 8206 11394 8258 11406
rect 8206 11330 8258 11342
rect 8542 11394 8594 11406
rect 8542 11330 8594 11342
rect 8766 11394 8818 11406
rect 8766 11330 8818 11342
rect 14366 11394 14418 11406
rect 31502 11394 31554 11406
rect 14802 11342 14814 11394
rect 14866 11342 14878 11394
rect 15810 11342 15822 11394
rect 15874 11342 15886 11394
rect 16930 11342 16942 11394
rect 16994 11342 17006 11394
rect 21522 11342 21534 11394
rect 21586 11342 21598 11394
rect 26002 11342 26014 11394
rect 26066 11342 26078 11394
rect 14366 11330 14418 11342
rect 31502 11330 31554 11342
rect 31726 11394 31778 11406
rect 42254 11394 42306 11406
rect 41906 11342 41918 11394
rect 41970 11342 41982 11394
rect 31726 11330 31778 11342
rect 42254 11330 42306 11342
rect 4958 11282 5010 11294
rect 4958 11218 5010 11230
rect 5070 11282 5122 11294
rect 5070 11218 5122 11230
rect 5630 11282 5682 11294
rect 5630 11218 5682 11230
rect 8654 11282 8706 11294
rect 8654 11218 8706 11230
rect 9214 11282 9266 11294
rect 9214 11218 9266 11230
rect 9326 11282 9378 11294
rect 9326 11218 9378 11230
rect 11006 11282 11058 11294
rect 11006 11218 11058 11230
rect 14030 11282 14082 11294
rect 14030 11218 14082 11230
rect 15150 11282 15202 11294
rect 31950 11282 32002 11294
rect 15362 11230 15374 11282
rect 15426 11230 15438 11282
rect 26226 11230 26238 11282
rect 26290 11230 26302 11282
rect 15150 11218 15202 11230
rect 31950 11218 32002 11230
rect 32174 11282 32226 11294
rect 32174 11218 32226 11230
rect 32398 11282 32450 11294
rect 32398 11218 32450 11230
rect 32510 11282 32562 11294
rect 32510 11218 32562 11230
rect 38222 11282 38274 11294
rect 38222 11218 38274 11230
rect 42590 11282 42642 11294
rect 52894 11282 52946 11294
rect 48850 11230 48862 11282
rect 48914 11230 48926 11282
rect 42590 11218 42642 11230
rect 52894 11218 52946 11230
rect 53230 11282 53282 11294
rect 53230 11218 53282 11230
rect 5742 11170 5794 11182
rect 5742 11106 5794 11118
rect 6974 11170 7026 11182
rect 6974 11106 7026 11118
rect 8990 11170 9042 11182
rect 8990 11106 9042 11118
rect 11342 11170 11394 11182
rect 11342 11106 11394 11118
rect 14142 11170 14194 11182
rect 14142 11106 14194 11118
rect 15262 11170 15314 11182
rect 15262 11106 15314 11118
rect 16606 11170 16658 11182
rect 16606 11106 16658 11118
rect 24782 11170 24834 11182
rect 24782 11106 24834 11118
rect 36206 11170 36258 11182
rect 36206 11106 36258 11118
rect 40798 11170 40850 11182
rect 40798 11106 40850 11118
rect 48526 11170 48578 11182
rect 48526 11106 48578 11118
rect 49982 11170 50034 11182
rect 49982 11106 50034 11118
rect 1344 11002 53648 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 50558 11002
rect 50610 10950 50662 11002
rect 50714 10950 50766 11002
rect 50818 10950 53648 11002
rect 1344 10916 53648 10950
rect 5070 10834 5122 10846
rect 5070 10770 5122 10782
rect 10894 10834 10946 10846
rect 10894 10770 10946 10782
rect 12014 10834 12066 10846
rect 12014 10770 12066 10782
rect 13246 10834 13298 10846
rect 13246 10770 13298 10782
rect 20750 10834 20802 10846
rect 20750 10770 20802 10782
rect 27358 10834 27410 10846
rect 27358 10770 27410 10782
rect 27918 10834 27970 10846
rect 27918 10770 27970 10782
rect 39454 10834 39506 10846
rect 39454 10770 39506 10782
rect 39902 10834 39954 10846
rect 39902 10770 39954 10782
rect 42702 10834 42754 10846
rect 42702 10770 42754 10782
rect 11678 10722 11730 10734
rect 2482 10670 2494 10722
rect 2546 10670 2558 10722
rect 11678 10658 11730 10670
rect 12798 10722 12850 10734
rect 12798 10658 12850 10670
rect 20974 10722 21026 10734
rect 27246 10722 27298 10734
rect 25218 10670 25230 10722
rect 25282 10670 25294 10722
rect 20974 10658 21026 10670
rect 27246 10658 27298 10670
rect 21086 10610 21138 10622
rect 1810 10558 1822 10610
rect 1874 10558 1886 10610
rect 10994 10558 11006 10610
rect 11058 10558 11070 10610
rect 11442 10558 11454 10610
rect 11506 10558 11518 10610
rect 12114 10558 12126 10610
rect 12178 10558 12190 10610
rect 12562 10558 12574 10610
rect 12626 10558 12638 10610
rect 21086 10546 21138 10558
rect 25566 10610 25618 10622
rect 25566 10546 25618 10558
rect 41022 10610 41074 10622
rect 41022 10546 41074 10558
rect 42814 10610 42866 10622
rect 42814 10546 42866 10558
rect 44270 10610 44322 10622
rect 44270 10546 44322 10558
rect 44494 10610 44546 10622
rect 45726 10610 45778 10622
rect 44818 10558 44830 10610
rect 44882 10558 44894 10610
rect 44494 10546 44546 10558
rect 45726 10546 45778 10558
rect 46398 10610 46450 10622
rect 47182 10610 47234 10622
rect 46610 10558 46622 10610
rect 46674 10558 46686 10610
rect 46398 10546 46450 10558
rect 47182 10546 47234 10558
rect 49198 10610 49250 10622
rect 49646 10610 49698 10622
rect 49410 10558 49422 10610
rect 49474 10558 49486 10610
rect 49746 10558 49758 10610
rect 49810 10558 49822 10610
rect 50306 10558 50318 10610
rect 50370 10558 50382 10610
rect 49198 10546 49250 10558
rect 49646 10546 49698 10558
rect 26014 10498 26066 10510
rect 4610 10446 4622 10498
rect 4674 10446 4686 10498
rect 26014 10434 26066 10446
rect 41582 10498 41634 10510
rect 41582 10434 41634 10446
rect 43262 10498 43314 10510
rect 43262 10434 43314 10446
rect 44382 10498 44434 10510
rect 48974 10498 49026 10510
rect 45266 10446 45278 10498
rect 45330 10446 45342 10498
rect 44382 10434 44434 10446
rect 48974 10434 49026 10446
rect 49310 10498 49362 10510
rect 51090 10446 51102 10498
rect 51154 10446 51166 10498
rect 53218 10446 53230 10498
rect 53282 10446 53294 10498
rect 49310 10434 49362 10446
rect 27358 10386 27410 10398
rect 42702 10386 42754 10398
rect 11106 10334 11118 10386
rect 11170 10334 11182 10386
rect 12226 10334 12238 10386
rect 12290 10334 12302 10386
rect 39218 10334 39230 10386
rect 39282 10383 39294 10386
rect 39890 10383 39902 10386
rect 39282 10337 39902 10383
rect 39282 10334 39294 10337
rect 39890 10334 39902 10337
rect 39954 10334 39966 10386
rect 27358 10322 27410 10334
rect 42702 10322 42754 10334
rect 1344 10218 53648 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 53648 10218
rect 1344 10132 53648 10166
rect 15934 10050 15986 10062
rect 15934 9986 15986 9998
rect 21422 10050 21474 10062
rect 21422 9986 21474 9998
rect 21982 10050 22034 10062
rect 21982 9986 22034 9998
rect 35422 10050 35474 10062
rect 35422 9986 35474 9998
rect 36206 10050 36258 10062
rect 50878 10050 50930 10062
rect 45042 9998 45054 10050
rect 45106 9998 45118 10050
rect 47058 9998 47070 10050
rect 47122 9998 47134 10050
rect 36206 9986 36258 9998
rect 50878 9986 50930 9998
rect 12014 9938 12066 9950
rect 7746 9886 7758 9938
rect 7810 9886 7822 9938
rect 9874 9886 9886 9938
rect 9938 9886 9950 9938
rect 12014 9874 12066 9886
rect 26462 9938 26514 9950
rect 50766 9938 50818 9950
rect 30258 9886 30270 9938
rect 30322 9886 30334 9938
rect 34850 9886 34862 9938
rect 34914 9886 34926 9938
rect 45154 9886 45166 9938
rect 45218 9886 45230 9938
rect 26462 9874 26514 9886
rect 50766 9874 50818 9886
rect 21310 9826 21362 9838
rect 6962 9774 6974 9826
rect 7026 9774 7038 9826
rect 21310 9762 21362 9774
rect 22094 9826 22146 9838
rect 22094 9762 22146 9774
rect 22766 9826 22818 9838
rect 22766 9762 22818 9774
rect 23102 9826 23154 9838
rect 27358 9826 27410 9838
rect 25778 9774 25790 9826
rect 25842 9774 25854 9826
rect 23102 9762 23154 9774
rect 27358 9762 27410 9774
rect 28030 9826 28082 9838
rect 28030 9762 28082 9774
rect 32734 9826 32786 9838
rect 32734 9762 32786 9774
rect 33406 9826 33458 9838
rect 33406 9762 33458 9774
rect 33854 9826 33906 9838
rect 33854 9762 33906 9774
rect 35646 9826 35698 9838
rect 38670 9826 38722 9838
rect 37090 9774 37102 9826
rect 37154 9774 37166 9826
rect 38210 9774 38222 9826
rect 38274 9774 38286 9826
rect 35646 9762 35698 9774
rect 38670 9762 38722 9774
rect 39006 9826 39058 9838
rect 39006 9762 39058 9774
rect 39230 9826 39282 9838
rect 45054 9826 45106 9838
rect 41458 9774 41470 9826
rect 41522 9774 41534 9826
rect 41906 9774 41918 9826
rect 41970 9774 41982 9826
rect 45490 9774 45502 9826
rect 45554 9774 45566 9826
rect 46834 9774 46846 9826
rect 46898 9774 46910 9826
rect 47394 9774 47406 9826
rect 47458 9774 47470 9826
rect 47954 9774 47966 9826
rect 48018 9774 48030 9826
rect 39230 9762 39282 9774
rect 45054 9762 45106 9774
rect 16046 9714 16098 9726
rect 16046 9650 16098 9662
rect 27806 9714 27858 9726
rect 27806 9650 27858 9662
rect 32958 9714 33010 9726
rect 32958 9650 33010 9662
rect 33518 9714 33570 9726
rect 33518 9650 33570 9662
rect 34638 9714 34690 9726
rect 34638 9650 34690 9662
rect 35982 9714 36034 9726
rect 40462 9714 40514 9726
rect 49198 9714 49250 9726
rect 49870 9714 49922 9726
rect 37986 9662 37998 9714
rect 38050 9662 38062 9714
rect 43586 9662 43598 9714
rect 43650 9662 43662 9714
rect 46946 9662 46958 9714
rect 47010 9662 47022 9714
rect 48850 9662 48862 9714
rect 48914 9662 48926 9714
rect 49522 9662 49534 9714
rect 49586 9662 49598 9714
rect 35982 9650 36034 9662
rect 40462 9650 40514 9662
rect 49198 9650 49250 9662
rect 49870 9650 49922 9662
rect 10334 9602 10386 9614
rect 10334 9538 10386 9550
rect 16718 9602 16770 9614
rect 16718 9538 16770 9550
rect 21422 9602 21474 9614
rect 21422 9538 21474 9550
rect 21982 9602 22034 9614
rect 21982 9538 22034 9550
rect 22878 9602 22930 9614
rect 27694 9602 27746 9614
rect 26002 9550 26014 9602
rect 26066 9550 26078 9602
rect 22878 9538 22930 9550
rect 27694 9538 27746 9550
rect 30718 9602 30770 9614
rect 30718 9538 30770 9550
rect 31166 9602 31218 9614
rect 31166 9538 31218 9550
rect 33070 9602 33122 9614
rect 33070 9538 33122 9550
rect 33742 9602 33794 9614
rect 33742 9538 33794 9550
rect 35310 9602 35362 9614
rect 38894 9602 38946 9614
rect 44270 9602 44322 9614
rect 37314 9550 37326 9602
rect 37378 9550 37390 9602
rect 40114 9550 40126 9602
rect 40178 9550 40190 9602
rect 35310 9538 35362 9550
rect 38894 9538 38946 9550
rect 44270 9538 44322 9550
rect 1344 9434 53648 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 50558 9434
rect 50610 9382 50662 9434
rect 50714 9382 50766 9434
rect 50818 9382 53648 9434
rect 1344 9348 53648 9382
rect 7310 9266 7362 9278
rect 7310 9202 7362 9214
rect 7758 9266 7810 9278
rect 7758 9202 7810 9214
rect 13246 9266 13298 9278
rect 13246 9202 13298 9214
rect 25342 9266 25394 9278
rect 25342 9202 25394 9214
rect 31502 9266 31554 9278
rect 31502 9202 31554 9214
rect 35646 9266 35698 9278
rect 35646 9202 35698 9214
rect 35870 9266 35922 9278
rect 35870 9202 35922 9214
rect 37662 9266 37714 9278
rect 46622 9266 46674 9278
rect 42690 9214 42702 9266
rect 42754 9214 42766 9266
rect 46162 9214 46174 9266
rect 46226 9214 46238 9266
rect 52882 9214 52894 9266
rect 52946 9214 52958 9266
rect 37662 9202 37714 9214
rect 46622 9202 46674 9214
rect 25566 9154 25618 9166
rect 35422 9154 35474 9166
rect 4722 9102 4734 9154
rect 4786 9102 4798 9154
rect 10658 9102 10670 9154
rect 10722 9102 10734 9154
rect 14354 9102 14366 9154
rect 14418 9102 14430 9154
rect 27682 9102 27694 9154
rect 27746 9102 27758 9154
rect 25566 9090 25618 9102
rect 35422 9090 35474 9102
rect 25678 9042 25730 9054
rect 39902 9042 39954 9054
rect 4050 8990 4062 9042
rect 4114 8990 4126 9042
rect 9874 8990 9886 9042
rect 9938 8990 9950 9042
rect 13682 8990 13694 9042
rect 13746 8990 13758 9042
rect 17378 8990 17390 9042
rect 17442 8990 17454 9042
rect 27010 8990 27022 9042
rect 27074 8990 27086 9042
rect 30930 8990 30942 9042
rect 30994 8990 31006 9042
rect 25678 8978 25730 8990
rect 39902 8978 39954 8990
rect 40350 9042 40402 9054
rect 43038 9042 43090 9054
rect 45726 9042 45778 9054
rect 53230 9042 53282 9054
rect 41682 8990 41694 9042
rect 41746 8990 41758 9042
rect 45490 8990 45502 9042
rect 45554 8990 45566 9042
rect 49410 8990 49422 9042
rect 49474 8990 49486 9042
rect 40350 8978 40402 8990
rect 43038 8978 43090 8990
rect 45726 8978 45778 8990
rect 53230 8978 53282 8990
rect 7198 8930 7250 8942
rect 13134 8930 13186 8942
rect 26574 8930 26626 8942
rect 30718 8930 30770 8942
rect 6850 8878 6862 8930
rect 6914 8878 6926 8930
rect 12786 8878 12798 8930
rect 12850 8878 12862 8930
rect 16482 8878 16494 8930
rect 16546 8878 16558 8930
rect 18162 8878 18174 8930
rect 18226 8878 18238 8930
rect 20290 8878 20302 8930
rect 20354 8878 20366 8930
rect 29810 8878 29822 8930
rect 29874 8878 29886 8930
rect 7198 8866 7250 8878
rect 13134 8866 13186 8878
rect 26574 8866 26626 8878
rect 30718 8866 30770 8878
rect 35534 8930 35586 8942
rect 48750 8930 48802 8942
rect 52670 8930 52722 8942
rect 41458 8878 41470 8930
rect 41522 8878 41534 8930
rect 45378 8878 45390 8930
rect 45442 8878 45454 8930
rect 49522 8878 49534 8930
rect 49586 8878 49598 8930
rect 35534 8866 35586 8878
rect 48750 8866 48802 8878
rect 52670 8866 52722 8878
rect 30606 8818 30658 8830
rect 39666 8766 39678 8818
rect 39730 8766 39742 8818
rect 41234 8766 41246 8818
rect 41298 8766 41310 8818
rect 30606 8754 30658 8766
rect 1344 8650 53648 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 53648 8650
rect 1344 8564 53648 8598
rect 13582 8370 13634 8382
rect 13582 8306 13634 8318
rect 17054 8370 17106 8382
rect 41470 8370 41522 8382
rect 45838 8370 45890 8382
rect 19394 8318 19406 8370
rect 19458 8318 19470 8370
rect 25890 8318 25902 8370
rect 25954 8318 25966 8370
rect 32386 8318 32398 8370
rect 32450 8318 32462 8370
rect 34514 8318 34526 8370
rect 34578 8318 34590 8370
rect 45378 8318 45390 8370
rect 45442 8318 45454 8370
rect 17054 8306 17106 8318
rect 41470 8306 41522 8318
rect 45838 8306 45890 8318
rect 49310 8370 49362 8382
rect 49310 8306 49362 8318
rect 7870 8258 7922 8270
rect 7870 8194 7922 8206
rect 8542 8258 8594 8270
rect 8542 8194 8594 8206
rect 8990 8258 9042 8270
rect 20526 8258 20578 8270
rect 22206 8258 22258 8270
rect 30494 8258 30546 8270
rect 20066 8206 20078 8258
rect 20130 8206 20142 8258
rect 20738 8206 20750 8258
rect 20802 8206 20814 8258
rect 22642 8206 22654 8258
rect 22706 8206 22718 8258
rect 23090 8206 23102 8258
rect 23154 8206 23166 8258
rect 8990 8194 9042 8206
rect 20526 8194 20578 8206
rect 22206 8194 22258 8206
rect 30494 8194 30546 8206
rect 31278 8258 31330 8270
rect 47742 8258 47794 8270
rect 49086 8258 49138 8270
rect 31602 8206 31614 8258
rect 31666 8206 31678 8258
rect 41010 8206 41022 8258
rect 41074 8206 41086 8258
rect 45154 8206 45166 8258
rect 45218 8206 45230 8258
rect 48850 8206 48862 8258
rect 48914 8206 48926 8258
rect 31278 8194 31330 8206
rect 47742 8194 47794 8206
rect 49086 8194 49138 8206
rect 8654 8146 8706 8158
rect 8654 8082 8706 8094
rect 8878 8146 8930 8158
rect 8878 8082 8930 8094
rect 19742 8146 19794 8158
rect 19742 8082 19794 8094
rect 20414 8146 20466 8158
rect 38334 8146 38386 8158
rect 23762 8094 23774 8146
rect 23826 8094 23838 8146
rect 20414 8082 20466 8094
rect 38334 8082 38386 8094
rect 41806 8146 41858 8158
rect 41806 8082 41858 8094
rect 41918 8146 41970 8158
rect 41918 8082 41970 8094
rect 48078 8146 48130 8158
rect 48078 8082 48130 8094
rect 48638 8146 48690 8158
rect 48638 8082 48690 8094
rect 49534 8146 49586 8158
rect 49534 8082 49586 8094
rect 50542 8146 50594 8158
rect 50542 8082 50594 8094
rect 7982 8034 8034 8046
rect 7982 7970 8034 7982
rect 8094 8034 8146 8046
rect 8094 7970 8146 7982
rect 9550 8034 9602 8046
rect 9550 7970 9602 7982
rect 19518 8034 19570 8046
rect 19518 7970 19570 7982
rect 20302 8034 20354 8046
rect 20302 7970 20354 7982
rect 22094 8034 22146 8046
rect 22094 7970 22146 7982
rect 22318 8034 22370 8046
rect 22318 7970 22370 7982
rect 22430 8034 22482 8046
rect 22430 7970 22482 7982
rect 26350 8034 26402 8046
rect 26350 7970 26402 7982
rect 30158 8034 30210 8046
rect 30158 7970 30210 7982
rect 37998 8034 38050 8046
rect 37998 7970 38050 7982
rect 38222 8034 38274 8046
rect 38222 7970 38274 7982
rect 42142 8034 42194 8046
rect 42142 7970 42194 7982
rect 42478 8034 42530 8046
rect 42478 7970 42530 7982
rect 48190 8034 48242 8046
rect 48190 7970 48242 7982
rect 48414 8034 48466 8046
rect 48414 7970 48466 7982
rect 49646 8034 49698 8046
rect 49646 7970 49698 7982
rect 50654 8034 50706 8046
rect 53006 8034 53058 8046
rect 52658 7982 52670 8034
rect 52722 7982 52734 8034
rect 50654 7970 50706 7982
rect 53006 7970 53058 7982
rect 1344 7866 53648 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 50558 7866
rect 50610 7814 50662 7866
rect 50714 7814 50766 7866
rect 50818 7814 53648 7866
rect 1344 7780 53648 7814
rect 8318 7698 8370 7710
rect 8318 7634 8370 7646
rect 8990 7698 9042 7710
rect 8990 7634 9042 7646
rect 13918 7698 13970 7710
rect 13918 7634 13970 7646
rect 20078 7698 20130 7710
rect 20078 7634 20130 7646
rect 20862 7698 20914 7710
rect 20862 7634 20914 7646
rect 23550 7698 23602 7710
rect 29374 7698 29426 7710
rect 33182 7698 33234 7710
rect 29026 7646 29038 7698
rect 29090 7646 29102 7698
rect 30258 7646 30270 7698
rect 30322 7646 30334 7698
rect 23550 7634 23602 7646
rect 29374 7634 29426 7646
rect 33182 7634 33234 7646
rect 35982 7698 36034 7710
rect 35982 7634 36034 7646
rect 41022 7698 41074 7710
rect 41022 7634 41074 7646
rect 42366 7698 42418 7710
rect 42366 7634 42418 7646
rect 43374 7698 43426 7710
rect 43374 7634 43426 7646
rect 44046 7698 44098 7710
rect 44046 7634 44098 7646
rect 44270 7698 44322 7710
rect 44270 7634 44322 7646
rect 48078 7698 48130 7710
rect 48078 7634 48130 7646
rect 48638 7698 48690 7710
rect 48638 7634 48690 7646
rect 8206 7586 8258 7598
rect 8206 7522 8258 7534
rect 19630 7586 19682 7598
rect 23326 7586 23378 7598
rect 27582 7586 27634 7598
rect 42142 7586 42194 7598
rect 21970 7534 21982 7586
rect 22034 7534 22046 7586
rect 27234 7534 27246 7586
rect 27298 7534 27310 7586
rect 39554 7534 39566 7586
rect 39618 7534 39630 7586
rect 19630 7522 19682 7534
rect 23326 7522 23378 7534
rect 27582 7522 27634 7534
rect 42142 7522 42194 7534
rect 42814 7586 42866 7598
rect 47742 7586 47794 7598
rect 45490 7534 45502 7586
rect 45554 7534 45566 7586
rect 46498 7534 46510 7586
rect 46562 7534 46574 7586
rect 42814 7522 42866 7534
rect 47742 7522 47794 7534
rect 47966 7586 48018 7598
rect 51090 7534 51102 7586
rect 51154 7534 51166 7586
rect 47966 7522 48018 7534
rect 8542 7474 8594 7486
rect 8542 7410 8594 7422
rect 19854 7474 19906 7486
rect 19854 7410 19906 7422
rect 20190 7474 20242 7486
rect 20190 7410 20242 7422
rect 22318 7474 22370 7486
rect 42590 7474 42642 7486
rect 48190 7474 48242 7486
rect 30034 7422 30046 7474
rect 30098 7422 30110 7474
rect 40338 7422 40350 7474
rect 40402 7422 40414 7474
rect 44818 7422 44830 7474
rect 44882 7422 44894 7474
rect 45714 7422 45726 7474
rect 45778 7422 45790 7474
rect 46274 7422 46286 7474
rect 46338 7422 46350 7474
rect 22318 7410 22370 7422
rect 42590 7410 42642 7422
rect 48190 7410 48242 7422
rect 49310 7474 49362 7486
rect 49310 7410 49362 7422
rect 49534 7474 49586 7486
rect 49534 7410 49586 7422
rect 49982 7474 50034 7486
rect 50306 7422 50318 7474
rect 50370 7422 50382 7474
rect 49982 7410 50034 7422
rect 14030 7362 14082 7374
rect 14030 7298 14082 7310
rect 19966 7362 20018 7374
rect 19966 7298 20018 7310
rect 20638 7362 20690 7374
rect 20638 7298 20690 7310
rect 20750 7362 20802 7374
rect 23650 7310 23662 7362
rect 23714 7310 23726 7362
rect 37426 7310 37438 7362
rect 37490 7310 37502 7362
rect 53218 7310 53230 7362
rect 53282 7310 53294 7362
rect 20750 7298 20802 7310
rect 42254 7250 42306 7262
rect 42254 7186 42306 7198
rect 49086 7250 49138 7262
rect 49086 7186 49138 7198
rect 1344 7082 53648 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 53648 7082
rect 1344 6996 53648 7030
rect 26798 6914 26850 6926
rect 26798 6850 26850 6862
rect 37550 6914 37602 6926
rect 37550 6850 37602 6862
rect 37774 6914 37826 6926
rect 37774 6850 37826 6862
rect 38222 6914 38274 6926
rect 38222 6850 38274 6862
rect 42254 6914 42306 6926
rect 42254 6850 42306 6862
rect 42926 6914 42978 6926
rect 42926 6850 42978 6862
rect 49870 6914 49922 6926
rect 49870 6850 49922 6862
rect 53006 6914 53058 6926
rect 53006 6850 53058 6862
rect 32174 6802 32226 6814
rect 36094 6802 36146 6814
rect 8530 6750 8542 6802
rect 8594 6750 8606 6802
rect 18274 6750 18286 6802
rect 18338 6750 18350 6802
rect 35746 6750 35758 6802
rect 35810 6750 35822 6802
rect 32174 6738 32226 6750
rect 36094 6738 36146 6750
rect 36206 6802 36258 6814
rect 36206 6738 36258 6750
rect 38334 6802 38386 6814
rect 38334 6738 38386 6750
rect 38782 6802 38834 6814
rect 38782 6738 38834 6750
rect 42030 6802 42082 6814
rect 50094 6802 50146 6814
rect 46050 6750 46062 6802
rect 46114 6750 46126 6802
rect 42030 6738 42082 6750
rect 50094 6738 50146 6750
rect 53230 6802 53282 6814
rect 53230 6738 53282 6750
rect 11342 6690 11394 6702
rect 7746 6638 7758 6690
rect 7810 6638 7822 6690
rect 11342 6626 11394 6638
rect 15038 6690 15090 6702
rect 27806 6690 27858 6702
rect 38222 6690 38274 6702
rect 15362 6638 15374 6690
rect 15426 6638 15438 6690
rect 16146 6638 16158 6690
rect 16210 6638 16222 6690
rect 25554 6638 25566 6690
rect 25618 6638 25630 6690
rect 29474 6638 29486 6690
rect 29538 6638 29550 6690
rect 32274 6638 32286 6690
rect 32338 6638 32350 6690
rect 32946 6638 32958 6690
rect 33010 6638 33022 6690
rect 36418 6638 36430 6690
rect 36482 6638 36494 6690
rect 15038 6626 15090 6638
rect 27806 6626 27858 6638
rect 38222 6626 38274 6638
rect 42478 6690 42530 6702
rect 49310 6690 49362 6702
rect 50318 6690 50370 6702
rect 46274 6638 46286 6690
rect 46338 6638 46350 6690
rect 49074 6638 49086 6690
rect 49138 6638 49150 6690
rect 49634 6638 49646 6690
rect 49698 6638 49710 6690
rect 42478 6626 42530 6638
rect 49310 6626 49362 6638
rect 50318 6626 50370 6638
rect 51550 6690 51602 6702
rect 51986 6638 51998 6690
rect 52050 6638 52062 6690
rect 51550 6626 51602 6638
rect 26910 6578 26962 6590
rect 25778 6526 25790 6578
rect 25842 6526 25854 6578
rect 26910 6514 26962 6526
rect 27470 6578 27522 6590
rect 27470 6514 27522 6526
rect 31726 6578 31778 6590
rect 39230 6578 39282 6590
rect 31938 6526 31950 6578
rect 32002 6526 32014 6578
rect 33618 6526 33630 6578
rect 33682 6526 33694 6578
rect 31726 6514 31778 6526
rect 39230 6514 39282 6526
rect 41806 6578 41858 6590
rect 45502 6578 45554 6590
rect 45154 6526 45166 6578
rect 45218 6526 45230 6578
rect 46722 6526 46734 6578
rect 46786 6526 46798 6578
rect 47394 6526 47406 6578
rect 47458 6526 47470 6578
rect 52658 6526 52670 6578
rect 52722 6526 52734 6578
rect 41806 6514 41858 6526
rect 45502 6514 45554 6526
rect 26798 6466 26850 6478
rect 10770 6414 10782 6466
rect 10834 6414 10846 6466
rect 26798 6402 26850 6414
rect 27582 6466 27634 6478
rect 32510 6466 32562 6478
rect 29250 6414 29262 6466
rect 29314 6414 29326 6466
rect 27582 6402 27634 6414
rect 32510 6402 32562 6414
rect 49870 6466 49922 6478
rect 49870 6402 49922 6414
rect 51326 6466 51378 6478
rect 51326 6402 51378 6414
rect 1344 6298 53648 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 50558 6298
rect 50610 6246 50662 6298
rect 50714 6246 50766 6298
rect 50818 6246 53648 6298
rect 1344 6212 53648 6246
rect 14702 6130 14754 6142
rect 14702 6066 14754 6078
rect 19742 6130 19794 6142
rect 19742 6066 19794 6078
rect 21646 6130 21698 6142
rect 21646 6066 21698 6078
rect 21758 6130 21810 6142
rect 21758 6066 21810 6078
rect 22430 6130 22482 6142
rect 22430 6066 22482 6078
rect 25566 6130 25618 6142
rect 25566 6066 25618 6078
rect 33070 6130 33122 6142
rect 33070 6066 33122 6078
rect 33294 6130 33346 6142
rect 33294 6066 33346 6078
rect 35870 6130 35922 6142
rect 35870 6066 35922 6078
rect 36878 6130 36930 6142
rect 36878 6066 36930 6078
rect 42702 6130 42754 6142
rect 42702 6066 42754 6078
rect 49198 6130 49250 6142
rect 49198 6066 49250 6078
rect 18958 6018 19010 6030
rect 12114 5966 12126 6018
rect 12178 5966 12190 6018
rect 18958 5954 19010 5966
rect 19966 6018 20018 6030
rect 19966 5954 20018 5966
rect 22878 6018 22930 6030
rect 36206 6018 36258 6030
rect 25218 5966 25230 6018
rect 25282 5966 25294 6018
rect 22878 5954 22930 5966
rect 36206 5954 36258 5966
rect 36318 6018 36370 6030
rect 36318 5954 36370 5966
rect 42030 6018 42082 6030
rect 42030 5954 42082 5966
rect 49870 6018 49922 6030
rect 49870 5954 49922 5966
rect 19630 5906 19682 5918
rect 21310 5906 21362 5918
rect 11330 5854 11342 5906
rect 11394 5854 11406 5906
rect 20178 5854 20190 5906
rect 20242 5854 20254 5906
rect 19630 5842 19682 5854
rect 21310 5842 21362 5854
rect 21422 5906 21474 5918
rect 22654 5906 22706 5918
rect 22194 5854 22206 5906
rect 22258 5854 22270 5906
rect 21422 5842 21474 5854
rect 22654 5842 22706 5854
rect 33742 5906 33794 5918
rect 33742 5842 33794 5854
rect 35982 5906 36034 5918
rect 35982 5842 36034 5854
rect 37214 5906 37266 5918
rect 37214 5842 37266 5854
rect 42366 5906 42418 5918
rect 42366 5842 42418 5854
rect 42590 5906 42642 5918
rect 50306 5854 50318 5906
rect 50370 5854 50382 5906
rect 42590 5842 42642 5854
rect 19854 5794 19906 5806
rect 14242 5742 14254 5794
rect 14306 5742 14318 5794
rect 19854 5730 19906 5742
rect 21534 5794 21586 5806
rect 21534 5730 21586 5742
rect 22542 5794 22594 5806
rect 22542 5730 22594 5742
rect 33182 5794 33234 5806
rect 33182 5730 33234 5742
rect 49534 5794 49586 5806
rect 51090 5742 51102 5794
rect 51154 5742 51166 5794
rect 53218 5742 53230 5794
rect 53282 5742 53294 5794
rect 49534 5730 49586 5742
rect 18846 5682 18898 5694
rect 18846 5618 18898 5630
rect 19182 5682 19234 5694
rect 19182 5618 19234 5630
rect 41806 5682 41858 5694
rect 41806 5618 41858 5630
rect 49982 5682 50034 5694
rect 49982 5618 50034 5630
rect 1344 5514 53648 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 53648 5514
rect 1344 5428 53648 5462
rect 19182 5346 19234 5358
rect 19182 5282 19234 5294
rect 22766 5346 22818 5358
rect 22766 5282 22818 5294
rect 31502 5346 31554 5358
rect 31502 5282 31554 5294
rect 38334 5346 38386 5358
rect 38334 5282 38386 5294
rect 45614 5346 45666 5358
rect 45614 5282 45666 5294
rect 29374 5234 29426 5246
rect 15250 5182 15262 5234
rect 15314 5182 15326 5234
rect 17378 5182 17390 5234
rect 17442 5182 17454 5234
rect 18834 5182 18846 5234
rect 18898 5182 18910 5234
rect 22418 5182 22430 5234
rect 22482 5182 22494 5234
rect 29374 5170 29426 5182
rect 29598 5234 29650 5246
rect 29598 5170 29650 5182
rect 30606 5234 30658 5246
rect 30606 5170 30658 5182
rect 36430 5234 36482 5246
rect 36430 5170 36482 5182
rect 40574 5234 40626 5246
rect 40574 5170 40626 5182
rect 44830 5234 44882 5246
rect 44830 5170 44882 5182
rect 46622 5234 46674 5246
rect 46622 5170 46674 5182
rect 47630 5234 47682 5246
rect 48178 5182 48190 5234
rect 48242 5182 48254 5234
rect 47630 5170 47682 5182
rect 17838 5122 17890 5134
rect 26126 5122 26178 5134
rect 28254 5122 28306 5134
rect 29710 5122 29762 5134
rect 14578 5070 14590 5122
rect 14642 5070 14654 5122
rect 25778 5070 25790 5122
rect 25842 5070 25854 5122
rect 27906 5070 27918 5122
rect 27970 5070 27982 5122
rect 28578 5070 28590 5122
rect 28642 5070 28654 5122
rect 17838 5058 17890 5070
rect 26126 5058 26178 5070
rect 28254 5058 28306 5070
rect 29710 5058 29762 5070
rect 30158 5122 30210 5134
rect 30158 5058 30210 5070
rect 31614 5122 31666 5134
rect 37998 5122 38050 5134
rect 46286 5122 46338 5134
rect 37202 5070 37214 5122
rect 37266 5070 37278 5122
rect 38770 5070 38782 5122
rect 38834 5070 38846 5122
rect 46050 5070 46062 5122
rect 46114 5070 46126 5122
rect 31614 5058 31666 5070
rect 37998 5058 38050 5070
rect 46286 5058 46338 5070
rect 48638 5122 48690 5134
rect 48638 5058 48690 5070
rect 49086 5122 49138 5134
rect 49086 5058 49138 5070
rect 18958 5010 19010 5022
rect 18958 4946 19010 4958
rect 22542 5010 22594 5022
rect 22542 4946 22594 4958
rect 28142 5010 28194 5022
rect 28142 4946 28194 4958
rect 28366 5010 28418 5022
rect 28366 4946 28418 4958
rect 29150 5010 29202 5022
rect 38882 4958 38894 5010
rect 38946 4958 38958 5010
rect 46498 4958 46510 5010
rect 46562 4958 46574 5010
rect 29150 4946 29202 4958
rect 24670 4898 24722 4910
rect 24670 4834 24722 4846
rect 26014 4898 26066 4910
rect 37438 4898 37490 4910
rect 29698 4846 29710 4898
rect 29762 4846 29774 4898
rect 26014 4834 26066 4846
rect 37438 4834 37490 4846
rect 39790 4898 39842 4910
rect 39790 4834 39842 4846
rect 44942 4898 44994 4910
rect 44942 4834 44994 4846
rect 1344 4730 53648 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 50558 4730
rect 50610 4678 50662 4730
rect 50714 4678 50766 4730
rect 50818 4678 53648 4730
rect 1344 4644 53648 4678
rect 16830 4562 16882 4574
rect 40238 4562 40290 4574
rect 36082 4510 36094 4562
rect 36146 4510 36158 4562
rect 16830 4498 16882 4510
rect 40238 4498 40290 4510
rect 14926 4450 14978 4462
rect 47854 4450 47906 4462
rect 18162 4398 18174 4450
rect 18226 4398 18238 4450
rect 22306 4398 22318 4450
rect 22370 4398 22382 4450
rect 26002 4398 26014 4450
rect 26066 4398 26078 4450
rect 30034 4398 30046 4450
rect 30098 4398 30110 4450
rect 33842 4398 33854 4450
rect 33906 4398 33918 4450
rect 37650 4398 37662 4450
rect 37714 4398 37726 4450
rect 41682 4398 41694 4450
rect 41746 4398 41758 4450
rect 44930 4398 44942 4450
rect 44994 4398 45006 4450
rect 14926 4386 14978 4398
rect 47854 4386 47906 4398
rect 48190 4450 48242 4462
rect 50866 4398 50878 4450
rect 50930 4398 50942 4450
rect 48190 4386 48242 4398
rect 47518 4338 47570 4350
rect 14354 4286 14366 4338
rect 14418 4286 14430 4338
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 21634 4286 21646 4338
rect 21698 4286 21710 4338
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 29250 4286 29262 4338
rect 29314 4286 29326 4338
rect 33058 4286 33070 4338
rect 33122 4286 33134 4338
rect 36978 4286 36990 4338
rect 37042 4286 37054 4338
rect 41010 4286 41022 4338
rect 41074 4286 41086 4338
rect 44258 4286 44270 4338
rect 44322 4286 44334 4338
rect 51650 4286 51662 4338
rect 51714 4286 51726 4338
rect 47518 4274 47570 4286
rect 3614 4226 3666 4238
rect 3614 4162 3666 4174
rect 3726 4226 3778 4238
rect 28814 4226 28866 4238
rect 20290 4174 20302 4226
rect 20354 4174 20366 4226
rect 24434 4174 24446 4226
rect 24498 4174 24510 4226
rect 28130 4174 28142 4226
rect 28194 4174 28206 4226
rect 32162 4174 32174 4226
rect 32226 4174 32238 4226
rect 39778 4174 39790 4226
rect 39842 4174 39854 4226
rect 43810 4174 43822 4226
rect 43874 4174 43886 4226
rect 47058 4174 47070 4226
rect 47122 4174 47134 4226
rect 48738 4174 48750 4226
rect 48802 4174 48814 4226
rect 3726 4162 3778 4174
rect 28814 4162 28866 4174
rect 12126 4114 12178 4126
rect 12126 4050 12178 4062
rect 1344 3946 53648 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 53648 3946
rect 1344 3860 53648 3894
rect 12462 3666 12514 3678
rect 12462 3602 12514 3614
rect 25006 3666 25058 3678
rect 25006 3602 25058 3614
rect 29038 3666 29090 3678
rect 29038 3602 29090 3614
rect 29822 3666 29874 3678
rect 29822 3602 29874 3614
rect 36990 3666 37042 3678
rect 50430 3666 50482 3678
rect 40226 3614 40238 3666
rect 40290 3614 40302 3666
rect 36990 3602 37042 3614
rect 50430 3602 50482 3614
rect 52670 3666 52722 3678
rect 52670 3602 52722 3614
rect 35534 3554 35586 3566
rect 46958 3554 47010 3566
rect 11890 3502 11902 3554
rect 11954 3502 11966 3554
rect 35970 3502 35982 3554
rect 36034 3502 36046 3554
rect 47618 3502 47630 3554
rect 47682 3502 47694 3554
rect 48514 3502 48526 3554
rect 48578 3502 48590 3554
rect 35534 3490 35586 3502
rect 46958 3490 47010 3502
rect 2718 3442 2770 3454
rect 2718 3378 2770 3390
rect 2942 3442 2994 3454
rect 2942 3378 2994 3390
rect 3278 3442 3330 3454
rect 39342 3442 39394 3454
rect 10098 3390 10110 3442
rect 10162 3390 10174 3442
rect 3278 3378 3330 3390
rect 39342 3378 39394 3390
rect 39790 3442 39842 3454
rect 39790 3378 39842 3390
rect 43150 3442 43202 3454
rect 43150 3378 43202 3390
rect 43598 3442 43650 3454
rect 52446 3442 52498 3454
rect 43922 3390 43934 3442
rect 43986 3390 43998 3442
rect 43598 3378 43650 3390
rect 52446 3378 52498 3390
rect 53230 3442 53282 3454
rect 53230 3378 53282 3390
rect 16942 3330 16994 3342
rect 16942 3266 16994 3278
rect 20862 3330 20914 3342
rect 20862 3266 20914 3278
rect 25342 3330 25394 3342
rect 47394 3278 47406 3330
rect 47458 3278 47470 3330
rect 25342 3266 25394 3278
rect 1344 3162 53648 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 50558 3162
rect 50610 3110 50662 3162
rect 50714 3110 50766 3162
rect 50818 3110 53648 3162
rect 1344 3076 53648 3110
<< via1 >>
rect 50430 51886 50482 51938
rect 51662 51886 51714 51938
rect 19838 51718 19890 51770
rect 19942 51718 19994 51770
rect 20046 51718 20098 51770
rect 50558 51718 50610 51770
rect 50662 51718 50714 51770
rect 50766 51718 50818 51770
rect 41246 51550 41298 51602
rect 41470 51550 41522 51602
rect 50542 51550 50594 51602
rect 41806 51438 41858 51490
rect 49982 51326 50034 51378
rect 50430 51326 50482 51378
rect 50654 51326 50706 51378
rect 51214 51326 51266 51378
rect 51438 51326 51490 51378
rect 51662 51326 51714 51378
rect 49758 51214 49810 51266
rect 51326 51214 51378 51266
rect 4478 50934 4530 50986
rect 4582 50934 4634 50986
rect 4686 50934 4738 50986
rect 35198 50934 35250 50986
rect 35302 50934 35354 50986
rect 35406 50934 35458 50986
rect 51102 50766 51154 50818
rect 18510 50654 18562 50706
rect 31054 50654 31106 50706
rect 40350 50654 40402 50706
rect 41246 50654 41298 50706
rect 48302 50654 48354 50706
rect 15710 50542 15762 50594
rect 24334 50542 24386 50594
rect 24782 50542 24834 50594
rect 27134 50542 27186 50594
rect 27694 50542 27746 50594
rect 33966 50542 34018 50594
rect 37438 50542 37490 50594
rect 44158 50542 44210 50594
rect 45502 50542 45554 50594
rect 51662 50542 51714 50594
rect 16382 50430 16434 50482
rect 23998 50430 24050 50482
rect 24110 50430 24162 50482
rect 24558 50430 24610 50482
rect 25006 50430 25058 50482
rect 25118 50430 25170 50482
rect 27358 50430 27410 50482
rect 27582 50430 27634 50482
rect 33182 50430 33234 50482
rect 38222 50430 38274 50482
rect 43374 50430 43426 50482
rect 44942 50430 44994 50482
rect 46174 50430 46226 50482
rect 18958 50318 19010 50370
rect 34414 50318 34466 50370
rect 37102 50318 37154 50370
rect 48750 50318 48802 50370
rect 19838 50150 19890 50202
rect 19942 50150 19994 50202
rect 20046 50150 20098 50202
rect 50558 50150 50610 50202
rect 50662 50150 50714 50202
rect 50766 50150 50818 50202
rect 17726 49982 17778 50034
rect 24110 49982 24162 50034
rect 27582 49982 27634 50034
rect 37774 49982 37826 50034
rect 38446 49982 38498 50034
rect 49646 49982 49698 50034
rect 18510 49870 18562 49922
rect 20750 49870 20802 49922
rect 26910 49870 26962 49922
rect 27358 49870 27410 49922
rect 28590 49870 28642 49922
rect 31054 49870 31106 49922
rect 31950 49870 32002 49922
rect 42030 49870 42082 49922
rect 51102 49870 51154 49922
rect 17390 49758 17442 49810
rect 17726 49758 17778 49810
rect 18062 49758 18114 49810
rect 18734 49758 18786 49810
rect 20078 49758 20130 49810
rect 25230 49758 25282 49810
rect 25454 49758 25506 49810
rect 25678 49758 25730 49810
rect 25790 49758 25842 49810
rect 26462 49758 26514 49810
rect 26686 49758 26738 49810
rect 27246 49758 27298 49810
rect 27918 49758 27970 49810
rect 31278 49758 31330 49810
rect 33966 49758 34018 49810
rect 37438 49758 37490 49810
rect 37550 49758 37602 49810
rect 37886 49758 37938 49810
rect 38670 49758 38722 49810
rect 48750 49758 48802 49810
rect 50318 49758 50370 49810
rect 19630 49646 19682 49698
rect 22878 49646 22930 49698
rect 23214 49646 23266 49698
rect 25566 49646 25618 49698
rect 26798 49646 26850 49698
rect 30718 49646 30770 49698
rect 31726 49646 31778 49698
rect 32062 49646 32114 49698
rect 34750 49646 34802 49698
rect 36878 49646 36930 49698
rect 37662 49646 37714 49698
rect 42142 49646 42194 49698
rect 48302 49646 48354 49698
rect 49198 49646 49250 49698
rect 49982 49646 50034 49698
rect 53230 49646 53282 49698
rect 23438 49534 23490 49586
rect 23662 49534 23714 49586
rect 38334 49534 38386 49586
rect 41806 49534 41858 49586
rect 48974 49534 49026 49586
rect 4478 49366 4530 49418
rect 4582 49366 4634 49418
rect 4686 49366 4738 49418
rect 35198 49366 35250 49418
rect 35302 49366 35354 49418
rect 35406 49366 35458 49418
rect 19294 49198 19346 49250
rect 27134 49198 27186 49250
rect 35086 49198 35138 49250
rect 35422 49198 35474 49250
rect 16382 49086 16434 49138
rect 27246 49086 27298 49138
rect 38334 49086 38386 49138
rect 41246 49086 41298 49138
rect 47070 49086 47122 49138
rect 51886 49086 51938 49138
rect 13582 48974 13634 49026
rect 18174 48974 18226 49026
rect 19630 48974 19682 49026
rect 19966 48974 20018 49026
rect 38222 48974 38274 49026
rect 38558 48974 38610 49026
rect 40910 48974 40962 49026
rect 41134 48974 41186 49026
rect 48750 48974 48802 49026
rect 48974 48974 49026 49026
rect 49198 48974 49250 49026
rect 49758 48974 49810 49026
rect 14254 48862 14306 48914
rect 18398 48862 18450 48914
rect 18510 48862 18562 48914
rect 20302 48862 20354 48914
rect 35198 48862 35250 48914
rect 37998 48862 38050 48914
rect 41358 48862 41410 48914
rect 41582 48862 41634 48914
rect 46734 48862 46786 48914
rect 47182 48862 47234 48914
rect 16830 48750 16882 48802
rect 19406 48750 19458 48802
rect 20190 48750 20242 48802
rect 30942 48750 30994 48802
rect 37102 48750 37154 48802
rect 38446 48750 38498 48802
rect 46398 48750 46450 48802
rect 46958 48750 47010 48802
rect 48302 48750 48354 48802
rect 19838 48582 19890 48634
rect 19942 48582 19994 48634
rect 20046 48582 20098 48634
rect 50558 48582 50610 48634
rect 50662 48582 50714 48634
rect 50766 48582 50818 48634
rect 21534 48414 21586 48466
rect 22206 48414 22258 48466
rect 25678 48414 25730 48466
rect 27022 48414 27074 48466
rect 27134 48414 27186 48466
rect 39790 48414 39842 48466
rect 42142 48414 42194 48466
rect 46846 48414 46898 48466
rect 49982 48414 50034 48466
rect 50206 48414 50258 48466
rect 20078 48302 20130 48354
rect 20414 48302 20466 48354
rect 20638 48302 20690 48354
rect 22094 48302 22146 48354
rect 22318 48302 22370 48354
rect 24558 48302 24610 48354
rect 25566 48302 25618 48354
rect 47070 48302 47122 48354
rect 48750 48302 48802 48354
rect 21086 48190 21138 48242
rect 21310 48190 21362 48242
rect 21646 48190 21698 48242
rect 22654 48190 22706 48242
rect 23102 48190 23154 48242
rect 23998 48190 24050 48242
rect 24446 48190 24498 48242
rect 25230 48190 25282 48242
rect 25790 48190 25842 48242
rect 26238 48190 26290 48242
rect 26462 48190 26514 48242
rect 26910 48190 26962 48242
rect 27582 48190 27634 48242
rect 31950 48190 32002 48242
rect 40126 48190 40178 48242
rect 42478 48190 42530 48242
rect 42926 48190 42978 48242
rect 46510 48190 46562 48242
rect 46846 48190 46898 48242
rect 49870 48190 49922 48242
rect 51102 48190 51154 48242
rect 19518 48078 19570 48130
rect 20750 48078 20802 48130
rect 21422 48078 21474 48130
rect 31614 48078 31666 48130
rect 41022 48078 41074 48130
rect 41806 48078 41858 48130
rect 43598 48078 43650 48130
rect 45726 48078 45778 48130
rect 46174 48078 46226 48130
rect 48190 48078 48242 48130
rect 49310 48078 49362 48130
rect 19742 47966 19794 48018
rect 24222 47966 24274 48018
rect 31950 47966 32002 48018
rect 48974 47966 49026 48018
rect 53006 47966 53058 48018
rect 4478 47798 4530 47850
rect 4582 47798 4634 47850
rect 4686 47798 4738 47850
rect 35198 47798 35250 47850
rect 35302 47798 35354 47850
rect 35406 47798 35458 47850
rect 26574 47630 26626 47682
rect 43038 47630 43090 47682
rect 51326 47630 51378 47682
rect 51550 47630 51602 47682
rect 24110 47518 24162 47570
rect 25342 47518 25394 47570
rect 32062 47518 32114 47570
rect 33182 47518 33234 47570
rect 35310 47518 35362 47570
rect 38558 47518 38610 47570
rect 49646 47518 49698 47570
rect 51102 47518 51154 47570
rect 14030 47406 14082 47458
rect 14590 47406 14642 47458
rect 19294 47406 19346 47458
rect 19630 47406 19682 47458
rect 25118 47406 25170 47458
rect 25678 47406 25730 47458
rect 26014 47406 26066 47458
rect 26350 47406 26402 47458
rect 27022 47406 27074 47458
rect 27134 47406 27186 47458
rect 28254 47406 28306 47458
rect 29150 47406 29202 47458
rect 32398 47406 32450 47458
rect 41582 47406 41634 47458
rect 49982 47406 50034 47458
rect 14142 47294 14194 47346
rect 19406 47294 19458 47346
rect 23774 47294 23826 47346
rect 24446 47294 24498 47346
rect 24782 47294 24834 47346
rect 25454 47294 25506 47346
rect 27246 47294 27298 47346
rect 27694 47294 27746 47346
rect 27918 47294 27970 47346
rect 28142 47294 28194 47346
rect 29934 47294 29986 47346
rect 41918 47294 41970 47346
rect 42254 47294 42306 47346
rect 42702 47294 42754 47346
rect 42926 47294 42978 47346
rect 48750 47294 48802 47346
rect 50430 47294 50482 47346
rect 50766 47294 50818 47346
rect 14254 47182 14306 47234
rect 18846 47182 18898 47234
rect 23998 47182 24050 47234
rect 26238 47182 26290 47234
rect 35758 47182 35810 47234
rect 41806 47182 41858 47234
rect 42030 47182 42082 47234
rect 46174 47182 46226 47234
rect 48862 47182 48914 47234
rect 49086 47182 49138 47234
rect 50990 47182 51042 47234
rect 51662 47182 51714 47234
rect 19838 47014 19890 47066
rect 19942 47014 19994 47066
rect 20046 47014 20098 47066
rect 50558 47014 50610 47066
rect 50662 47014 50714 47066
rect 50766 47014 50818 47066
rect 13246 46846 13298 46898
rect 14702 46846 14754 46898
rect 21086 46846 21138 46898
rect 27470 46846 27522 46898
rect 27694 46846 27746 46898
rect 32286 46846 32338 46898
rect 38670 46846 38722 46898
rect 40014 46846 40066 46898
rect 12014 46734 12066 46786
rect 12238 46734 12290 46786
rect 14030 46734 14082 46786
rect 20078 46734 20130 46786
rect 20414 46734 20466 46786
rect 20974 46734 21026 46786
rect 23438 46734 23490 46786
rect 27358 46734 27410 46786
rect 30270 46734 30322 46786
rect 30942 46734 30994 46786
rect 33518 46734 33570 46786
rect 51102 46734 51154 46786
rect 12350 46622 12402 46674
rect 13134 46622 13186 46674
rect 13358 46622 13410 46674
rect 13806 46622 13858 46674
rect 14254 46622 14306 46674
rect 14478 46622 14530 46674
rect 14702 46622 14754 46674
rect 15038 46622 15090 46674
rect 18958 46622 19010 46674
rect 19630 46622 19682 46674
rect 20302 46622 20354 46674
rect 22542 46622 22594 46674
rect 24670 46622 24722 46674
rect 30158 46622 30210 46674
rect 33742 46622 33794 46674
rect 35534 46622 35586 46674
rect 38894 46622 38946 46674
rect 39342 46622 39394 46674
rect 40238 46622 40290 46674
rect 47182 46622 47234 46674
rect 48190 46622 48242 46674
rect 48750 46622 48802 46674
rect 50318 46622 50370 46674
rect 11902 46510 11954 46562
rect 12798 46510 12850 46562
rect 15150 46510 15202 46562
rect 29934 46510 29986 46562
rect 36206 46510 36258 46562
rect 38334 46510 38386 46562
rect 38782 46510 38834 46562
rect 39678 46510 39730 46562
rect 44382 46510 44434 46562
rect 46510 46510 46562 46562
rect 47742 46510 47794 46562
rect 49310 46510 49362 46562
rect 49982 46510 50034 46562
rect 53230 46510 53282 46562
rect 4478 46230 4530 46282
rect 4582 46230 4634 46282
rect 4686 46230 4738 46282
rect 35198 46230 35250 46282
rect 35302 46230 35354 46282
rect 35406 46230 35458 46282
rect 18958 46062 19010 46114
rect 19294 46062 19346 46114
rect 21870 46062 21922 46114
rect 44158 46062 44210 46114
rect 11566 45950 11618 46002
rect 14254 45950 14306 46002
rect 18734 45950 18786 46002
rect 22542 45950 22594 46002
rect 37102 45950 37154 46002
rect 38558 45950 38610 46002
rect 42366 45950 42418 46002
rect 8766 45838 8818 45890
rect 12014 45838 12066 45890
rect 14030 45838 14082 45890
rect 15038 45838 15090 45890
rect 15934 45838 15986 45890
rect 22430 45838 22482 45890
rect 22654 45838 22706 45890
rect 33966 45838 34018 45890
rect 34302 45838 34354 45890
rect 37550 45838 37602 45890
rect 38222 45838 38274 45890
rect 39790 45838 39842 45890
rect 42030 45838 42082 45890
rect 43038 45838 43090 45890
rect 43262 45838 43314 45890
rect 43374 45838 43426 45890
rect 9438 45726 9490 45778
rect 14478 45726 14530 45778
rect 16606 45726 16658 45778
rect 24334 45726 24386 45778
rect 25006 45726 25058 45778
rect 36990 45726 37042 45778
rect 37326 45726 37378 45778
rect 37886 45726 37938 45778
rect 37998 45726 38050 45778
rect 39566 45726 39618 45778
rect 40574 45726 40626 45778
rect 41806 45726 41858 45778
rect 42366 45726 42418 45778
rect 43150 45726 43202 45778
rect 43822 45726 43874 45778
rect 49086 45726 49138 45778
rect 12126 45614 12178 45666
rect 12238 45614 12290 45666
rect 12462 45614 12514 45666
rect 13582 45614 13634 45666
rect 19182 45614 19234 45666
rect 23998 45614 24050 45666
rect 24670 45614 24722 45666
rect 25454 45614 25506 45666
rect 34078 45614 34130 45666
rect 40238 45614 40290 45666
rect 42254 45614 42306 45666
rect 42926 45614 42978 45666
rect 44046 45614 44098 45666
rect 49198 45614 49250 45666
rect 19838 45446 19890 45498
rect 19942 45446 19994 45498
rect 20046 45446 20098 45498
rect 50558 45446 50610 45498
rect 50662 45446 50714 45498
rect 50766 45446 50818 45498
rect 11566 45278 11618 45330
rect 12462 45278 12514 45330
rect 22878 45278 22930 45330
rect 23214 45278 23266 45330
rect 36542 45278 36594 45330
rect 37326 45278 37378 45330
rect 37998 45278 38050 45330
rect 41134 45278 41186 45330
rect 43150 45278 43202 45330
rect 49982 45278 50034 45330
rect 11790 45166 11842 45218
rect 14254 45166 14306 45218
rect 14366 45166 14418 45218
rect 18062 45166 18114 45218
rect 18622 45166 18674 45218
rect 19070 45166 19122 45218
rect 33406 45166 33458 45218
rect 33630 45166 33682 45218
rect 38334 45166 38386 45218
rect 38894 45166 38946 45218
rect 39454 45166 39506 45218
rect 42926 45166 42978 45218
rect 48190 45166 48242 45218
rect 50094 45166 50146 45218
rect 11342 45054 11394 45106
rect 11566 45054 11618 45106
rect 12238 45054 12290 45106
rect 14030 45054 14082 45106
rect 18286 45054 18338 45106
rect 18958 45054 19010 45106
rect 22654 45054 22706 45106
rect 23438 45054 23490 45106
rect 26014 45054 26066 45106
rect 32062 45054 32114 45106
rect 32286 45054 32338 45106
rect 34638 45054 34690 45106
rect 35422 45054 35474 45106
rect 35646 45054 35698 45106
rect 35758 45054 35810 45106
rect 37102 45054 37154 45106
rect 37438 45054 37490 45106
rect 38446 45054 38498 45106
rect 38782 45054 38834 45106
rect 40910 45054 40962 45106
rect 41358 45054 41410 45106
rect 41470 45054 41522 45106
rect 43822 45054 43874 45106
rect 47854 45054 47906 45106
rect 48974 45054 49026 45106
rect 49198 45054 49250 45106
rect 49758 45054 49810 45106
rect 51102 45054 51154 45106
rect 15374 44942 15426 44994
rect 18174 44942 18226 44994
rect 19742 44942 19794 44994
rect 24558 44942 24610 44994
rect 31502 44942 31554 44994
rect 34190 44942 34242 44994
rect 41246 44942 41298 44994
rect 43262 44942 43314 44994
rect 44494 44942 44546 44994
rect 46622 44942 46674 44994
rect 47070 44942 47122 44994
rect 47518 44942 47570 44994
rect 48078 44942 48130 44994
rect 48750 44942 48802 44994
rect 14814 44830 14866 44882
rect 19070 44830 19122 44882
rect 26126 44830 26178 44882
rect 33294 44830 33346 44882
rect 34302 44830 34354 44882
rect 36206 44830 36258 44882
rect 36430 44830 36482 44882
rect 53006 44830 53058 44882
rect 4478 44662 4530 44714
rect 4582 44662 4634 44714
rect 4686 44662 4738 44714
rect 35198 44662 35250 44714
rect 35302 44662 35354 44714
rect 35406 44662 35458 44714
rect 17278 44494 17330 44546
rect 17614 44494 17666 44546
rect 22094 44494 22146 44546
rect 26910 44494 26962 44546
rect 17726 44382 17778 44434
rect 18622 44382 18674 44434
rect 19406 44382 19458 44434
rect 26126 44382 26178 44434
rect 32062 44382 32114 44434
rect 32510 44382 32562 44434
rect 32846 44382 32898 44434
rect 33966 44382 34018 44434
rect 48526 44382 48578 44434
rect 16158 44270 16210 44322
rect 16830 44270 16882 44322
rect 17390 44270 17442 44322
rect 18174 44270 18226 44322
rect 18846 44270 18898 44322
rect 19854 44270 19906 44322
rect 20078 44270 20130 44322
rect 22206 44270 22258 44322
rect 22878 44270 22930 44322
rect 23438 44270 23490 44322
rect 25454 44270 25506 44322
rect 25790 44270 25842 44322
rect 29150 44270 29202 44322
rect 34750 44270 34802 44322
rect 35758 44270 35810 44322
rect 48974 44270 49026 44322
rect 16382 44158 16434 44210
rect 18398 44158 18450 44210
rect 22542 44158 22594 44210
rect 25118 44158 25170 44210
rect 29934 44158 29986 44210
rect 34862 44158 34914 44210
rect 36430 44158 36482 44210
rect 49422 44158 49474 44210
rect 50542 44158 50594 44210
rect 11566 44046 11618 44098
rect 19518 44046 19570 44098
rect 19966 44046 20018 44098
rect 20302 44046 20354 44098
rect 22094 44046 22146 44098
rect 23214 44046 23266 44098
rect 25454 44046 25506 44098
rect 26014 44046 26066 44098
rect 26238 44046 26290 44098
rect 26462 44046 26514 44098
rect 27022 44046 27074 44098
rect 27134 44046 27186 44098
rect 32958 44046 33010 44098
rect 33406 44046 33458 44098
rect 36318 44046 36370 44098
rect 38670 44046 38722 44098
rect 49982 44046 50034 44098
rect 50878 44046 50930 44098
rect 19838 43878 19890 43930
rect 19942 43878 19994 43930
rect 20046 43878 20098 43930
rect 50558 43878 50610 43930
rect 50662 43878 50714 43930
rect 50766 43878 50818 43930
rect 11230 43710 11282 43762
rect 18062 43710 18114 43762
rect 20190 43710 20242 43762
rect 21422 43710 21474 43762
rect 26126 43710 26178 43762
rect 29374 43710 29426 43762
rect 33742 43710 33794 43762
rect 34414 43710 34466 43762
rect 38894 43710 38946 43762
rect 46062 43710 46114 43762
rect 11790 43598 11842 43650
rect 12350 43598 12402 43650
rect 12574 43598 12626 43650
rect 14030 43598 14082 43650
rect 14142 43598 14194 43650
rect 18734 43598 18786 43650
rect 20078 43598 20130 43650
rect 20750 43598 20802 43650
rect 21086 43598 21138 43650
rect 26798 43598 26850 43650
rect 27918 43598 27970 43650
rect 28590 43598 28642 43650
rect 49646 43598 49698 43650
rect 51102 43598 51154 43650
rect 10894 43486 10946 43538
rect 11566 43486 11618 43538
rect 12238 43486 12290 43538
rect 12686 43486 12738 43538
rect 14366 43486 14418 43538
rect 14702 43486 14754 43538
rect 18286 43486 18338 43538
rect 18958 43486 19010 43538
rect 20414 43486 20466 43538
rect 25566 43486 25618 43538
rect 25902 43486 25954 43538
rect 27134 43486 27186 43538
rect 27358 43486 27410 43538
rect 28366 43486 28418 43538
rect 29262 43486 29314 43538
rect 33518 43486 33570 43538
rect 34078 43486 34130 43538
rect 38782 43486 38834 43538
rect 39118 43486 39170 43538
rect 45950 43486 46002 43538
rect 46286 43486 46338 43538
rect 49086 43486 49138 43538
rect 49310 43486 49362 43538
rect 50318 43486 50370 43538
rect 12014 43374 12066 43426
rect 18510 43374 18562 43426
rect 19854 43374 19906 43426
rect 25790 43374 25842 43426
rect 27246 43374 27298 43426
rect 34862 43374 34914 43426
rect 48302 43374 48354 43426
rect 53230 43374 53282 43426
rect 29038 43262 29090 43314
rect 29374 43262 29426 43314
rect 4478 43094 4530 43146
rect 4582 43094 4634 43146
rect 4686 43094 4738 43146
rect 35198 43094 35250 43146
rect 35302 43094 35354 43146
rect 35406 43094 35458 43146
rect 14030 42926 14082 42978
rect 14366 42926 14418 42978
rect 15262 42926 15314 42978
rect 29710 42926 29762 42978
rect 33966 42926 34018 42978
rect 38670 42926 38722 42978
rect 9662 42814 9714 42866
rect 11790 42814 11842 42866
rect 12238 42814 12290 42866
rect 16046 42814 16098 42866
rect 23662 42814 23714 42866
rect 43150 42814 43202 42866
rect 8878 42702 8930 42754
rect 14702 42702 14754 42754
rect 15374 42702 15426 42754
rect 24110 42702 24162 42754
rect 33070 42702 33122 42754
rect 33294 42702 33346 42754
rect 33518 42702 33570 42754
rect 36990 42702 37042 42754
rect 37774 42702 37826 42754
rect 38446 42702 38498 42754
rect 40350 42702 40402 42754
rect 44270 42702 44322 42754
rect 44830 42702 44882 42754
rect 45390 42702 45442 42754
rect 13806 42590 13858 42642
rect 14926 42590 14978 42642
rect 37102 42590 37154 42642
rect 37662 42590 37714 42642
rect 39006 42590 39058 42642
rect 39342 42590 39394 42642
rect 39678 42590 39730 42642
rect 41022 42590 41074 42642
rect 43486 42590 43538 42642
rect 45502 42590 45554 42642
rect 15150 42478 15202 42530
rect 23550 42478 23602 42530
rect 23774 42478 23826 42530
rect 28590 42478 28642 42530
rect 29822 42478 29874 42530
rect 29934 42478 29986 42530
rect 30494 42478 30546 42530
rect 32286 42478 32338 42530
rect 32734 42478 32786 42530
rect 37326 42478 37378 42530
rect 37438 42478 37490 42530
rect 43822 42478 43874 42530
rect 44942 42478 44994 42530
rect 45166 42478 45218 42530
rect 45726 42478 45778 42530
rect 49982 42478 50034 42530
rect 19838 42310 19890 42362
rect 19942 42310 19994 42362
rect 20046 42310 20098 42362
rect 50558 42310 50610 42362
rect 50662 42310 50714 42362
rect 50766 42310 50818 42362
rect 12686 42142 12738 42194
rect 14142 42142 14194 42194
rect 14366 42142 14418 42194
rect 15038 42142 15090 42194
rect 23550 42142 23602 42194
rect 27022 42142 27074 42194
rect 33182 42142 33234 42194
rect 38446 42142 38498 42194
rect 40014 42142 40066 42194
rect 41134 42142 41186 42194
rect 43262 42142 43314 42194
rect 49870 42142 49922 42194
rect 14590 42030 14642 42082
rect 15150 42030 15202 42082
rect 29822 42030 29874 42082
rect 38334 42030 38386 42082
rect 39902 42030 39954 42082
rect 43374 42030 43426 42082
rect 5070 41918 5122 41970
rect 12350 41918 12402 41970
rect 22990 41918 23042 41970
rect 23326 41918 23378 41970
rect 23774 41918 23826 41970
rect 23886 41918 23938 41970
rect 26126 41918 26178 41970
rect 26350 41918 26402 41970
rect 26798 41918 26850 41970
rect 27358 41918 27410 41970
rect 29150 41918 29202 41970
rect 33518 41918 33570 41970
rect 38670 41918 38722 41970
rect 40238 41918 40290 41970
rect 40910 41918 40962 41970
rect 41246 41918 41298 41970
rect 48078 41918 48130 41970
rect 48862 41918 48914 41970
rect 49310 41918 49362 41970
rect 50430 41918 50482 41970
rect 5742 41806 5794 41858
rect 7870 41806 7922 41858
rect 8318 41806 8370 41858
rect 23662 41806 23714 41858
rect 24446 41806 24498 41858
rect 26574 41806 26626 41858
rect 31950 41806 32002 41858
rect 36654 41806 36706 41858
rect 45278 41806 45330 41858
rect 47406 41806 47458 41858
rect 49870 41806 49922 41858
rect 51102 41806 51154 41858
rect 53230 41806 53282 41858
rect 14478 41694 14530 41746
rect 15038 41694 15090 41746
rect 22654 41694 22706 41746
rect 23102 41694 23154 41746
rect 24334 41694 24386 41746
rect 33182 41694 33234 41746
rect 33294 41694 33346 41746
rect 43262 41694 43314 41746
rect 49646 41694 49698 41746
rect 4478 41526 4530 41578
rect 4582 41526 4634 41578
rect 4686 41526 4738 41578
rect 35198 41526 35250 41578
rect 35302 41526 35354 41578
rect 35406 41526 35458 41578
rect 14814 41358 14866 41410
rect 26462 41358 26514 41410
rect 26798 41358 26850 41410
rect 17054 41246 17106 41298
rect 19182 41246 19234 41298
rect 24782 41246 24834 41298
rect 32398 41246 32450 41298
rect 36430 41246 36482 41298
rect 49086 41246 49138 41298
rect 51886 41246 51938 41298
rect 14366 41134 14418 41186
rect 14702 41134 14754 41186
rect 15150 41134 15202 41186
rect 16382 41134 16434 41186
rect 22206 41134 22258 41186
rect 22766 41134 22818 41186
rect 26014 41134 26066 41186
rect 26574 41134 26626 41186
rect 33518 41134 33570 41186
rect 37326 41134 37378 41186
rect 45614 41134 45666 41186
rect 48526 41134 48578 41186
rect 49198 41134 49250 41186
rect 49982 41134 50034 41186
rect 23438 41022 23490 41074
rect 24558 41022 24610 41074
rect 34302 41022 34354 41074
rect 36990 41022 37042 41074
rect 37102 41022 37154 41074
rect 37550 41022 37602 41074
rect 45278 41022 45330 41074
rect 45838 41022 45890 41074
rect 14478 40910 14530 40962
rect 15598 40910 15650 40962
rect 19630 40910 19682 40962
rect 22430 40910 22482 40962
rect 26462 40910 26514 40962
rect 27358 40910 27410 40962
rect 40574 40910 40626 40962
rect 41806 40910 41858 40962
rect 45726 40910 45778 40962
rect 48414 40910 48466 40962
rect 48974 40910 49026 40962
rect 19838 40742 19890 40794
rect 19942 40742 19994 40794
rect 20046 40742 20098 40794
rect 50558 40742 50610 40794
rect 50662 40742 50714 40794
rect 50766 40742 50818 40794
rect 5742 40574 5794 40626
rect 15374 40574 15426 40626
rect 22654 40574 22706 40626
rect 23326 40574 23378 40626
rect 24334 40574 24386 40626
rect 38894 40574 38946 40626
rect 42030 40574 42082 40626
rect 44046 40574 44098 40626
rect 44270 40574 44322 40626
rect 7982 40462 8034 40514
rect 19742 40462 19794 40514
rect 22990 40462 23042 40514
rect 23886 40462 23938 40514
rect 24222 40462 24274 40514
rect 26574 40462 26626 40514
rect 35310 40462 35362 40514
rect 38558 40462 38610 40514
rect 40126 40462 40178 40514
rect 41470 40462 41522 40514
rect 42366 40462 42418 40514
rect 43710 40462 43762 40514
rect 5406 40350 5458 40402
rect 5742 40350 5794 40402
rect 5966 40350 6018 40402
rect 8318 40350 8370 40402
rect 16606 40350 16658 40402
rect 18622 40350 18674 40402
rect 19070 40350 19122 40402
rect 23326 40350 23378 40402
rect 23438 40350 23490 40402
rect 23662 40350 23714 40402
rect 24558 40350 24610 40402
rect 25902 40350 25954 40402
rect 29150 40350 29202 40402
rect 31950 40350 32002 40402
rect 32174 40350 32226 40402
rect 33294 40350 33346 40402
rect 38110 40350 38162 40402
rect 40014 40350 40066 40402
rect 40798 40350 40850 40402
rect 41134 40350 41186 40402
rect 43934 40350 43986 40402
rect 44494 40350 44546 40402
rect 50654 40350 50706 40402
rect 15486 40238 15538 40290
rect 21870 40238 21922 40290
rect 28702 40238 28754 40290
rect 32398 40238 32450 40290
rect 35758 40238 35810 40290
rect 41022 40238 41074 40290
rect 46846 40238 46898 40290
rect 40126 40126 40178 40178
rect 53006 40126 53058 40178
rect 4478 39958 4530 40010
rect 4582 39958 4634 40010
rect 4686 39958 4738 40010
rect 35198 39958 35250 40010
rect 35302 39958 35354 40010
rect 35406 39958 35458 40010
rect 5966 39790 6018 39842
rect 6526 39790 6578 39842
rect 8430 39790 8482 39842
rect 37102 39790 37154 39842
rect 12798 39678 12850 39730
rect 14254 39678 14306 39730
rect 16382 39678 16434 39730
rect 17390 39678 17442 39730
rect 23998 39678 24050 39730
rect 27918 39678 27970 39730
rect 38446 39678 38498 39730
rect 40574 39678 40626 39730
rect 46734 39678 46786 39730
rect 9326 39566 9378 39618
rect 9550 39566 9602 39618
rect 9886 39566 9938 39618
rect 13582 39566 13634 39618
rect 17054 39566 17106 39618
rect 18958 39566 19010 39618
rect 19294 39566 19346 39618
rect 28366 39566 28418 39618
rect 41358 39566 41410 39618
rect 41806 39566 41858 39618
rect 44046 39566 44098 39618
rect 44718 39566 44770 39618
rect 45166 39566 45218 39618
rect 49646 39566 49698 39618
rect 50318 39566 50370 39618
rect 50766 39566 50818 39618
rect 50878 39566 50930 39618
rect 51326 39566 51378 39618
rect 4958 39454 5010 39506
rect 5630 39454 5682 39506
rect 6078 39454 6130 39506
rect 6414 39454 6466 39506
rect 6526 39454 6578 39506
rect 8094 39454 8146 39506
rect 8542 39454 8594 39506
rect 8990 39454 9042 39506
rect 9438 39454 9490 39506
rect 10670 39454 10722 39506
rect 17726 39454 17778 39506
rect 19406 39454 19458 39506
rect 36206 39454 36258 39506
rect 37102 39454 37154 39506
rect 37214 39454 37266 39506
rect 45390 39454 45442 39506
rect 46062 39454 46114 39506
rect 48862 39454 48914 39506
rect 52110 39454 52162 39506
rect 5070 39342 5122 39394
rect 5854 39342 5906 39394
rect 8318 39342 8370 39394
rect 36318 39342 36370 39394
rect 36542 39342 36594 39394
rect 44158 39342 44210 39394
rect 44382 39342 44434 39394
rect 44942 39342 44994 39394
rect 46174 39342 46226 39394
rect 46398 39342 46450 39394
rect 50206 39342 50258 39394
rect 50990 39342 51042 39394
rect 51438 39342 51490 39394
rect 51550 39342 51602 39394
rect 19838 39174 19890 39226
rect 19942 39174 19994 39226
rect 20046 39174 20098 39226
rect 50558 39174 50610 39226
rect 50662 39174 50714 39226
rect 50766 39174 50818 39226
rect 7198 39006 7250 39058
rect 9886 39006 9938 39058
rect 10110 39006 10162 39058
rect 13022 39006 13074 39058
rect 19518 39006 19570 39058
rect 34862 39006 34914 39058
rect 46398 39006 46450 39058
rect 46958 39006 47010 39058
rect 7982 38894 8034 38946
rect 8094 38894 8146 38946
rect 19742 38894 19794 38946
rect 22318 38894 22370 38946
rect 30942 38894 30994 38946
rect 32398 38894 32450 38946
rect 44942 38894 44994 38946
rect 47070 38894 47122 38946
rect 47294 38894 47346 38946
rect 51102 38894 51154 38946
rect 7534 38782 7586 38834
rect 8206 38782 8258 38834
rect 9774 38782 9826 38834
rect 16382 38782 16434 38834
rect 16606 38782 16658 38834
rect 17950 38782 18002 38834
rect 19854 38782 19906 38834
rect 20862 38782 20914 38834
rect 21646 38782 21698 38834
rect 30046 38782 30098 38834
rect 30494 38782 30546 38834
rect 30830 38782 30882 38834
rect 32510 38782 32562 38834
rect 33294 38782 33346 38834
rect 33742 38782 33794 38834
rect 37774 38782 37826 38834
rect 45726 38782 45778 38834
rect 46622 38782 46674 38834
rect 50430 38782 50482 38834
rect 16830 38670 16882 38722
rect 17390 38670 17442 38722
rect 8654 38558 8706 38610
rect 17614 38670 17666 38722
rect 20190 38670 20242 38722
rect 21086 38670 21138 38722
rect 24446 38670 24498 38722
rect 29262 38670 29314 38722
rect 29598 38670 29650 38722
rect 32062 38670 32114 38722
rect 33630 38670 33682 38722
rect 36318 38670 36370 38722
rect 42814 38670 42866 38722
rect 53230 38670 53282 38722
rect 17950 38558 18002 38610
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 5966 38222 6018 38274
rect 8766 38222 8818 38274
rect 17950 38222 18002 38274
rect 8542 38110 8594 38162
rect 19966 38110 20018 38162
rect 31390 38110 31442 38162
rect 36430 38110 36482 38162
rect 44270 38110 44322 38162
rect 45950 38110 46002 38162
rect 6078 37998 6130 38050
rect 18062 37998 18114 38050
rect 18286 37998 18338 38050
rect 18510 37998 18562 38050
rect 18622 37998 18674 38050
rect 19630 37998 19682 38050
rect 20190 37998 20242 38050
rect 25790 37998 25842 38050
rect 26350 37998 26402 38050
rect 28142 37998 28194 38050
rect 28478 37998 28530 38050
rect 30046 37998 30098 38050
rect 30494 37998 30546 38050
rect 30718 37998 30770 38050
rect 32286 37998 32338 38050
rect 33630 37998 33682 38050
rect 36990 37998 37042 38050
rect 37326 37998 37378 38050
rect 37550 37998 37602 38050
rect 44830 37998 44882 38050
rect 4958 37886 5010 37938
rect 5070 37886 5122 37938
rect 5966 37886 6018 37938
rect 9550 37886 9602 37938
rect 9662 37886 9714 37938
rect 19070 37886 19122 37938
rect 20638 37886 20690 37938
rect 26462 37886 26514 37938
rect 28590 37886 28642 37938
rect 31950 37886 32002 37938
rect 32062 37886 32114 37938
rect 34302 37886 34354 37938
rect 37102 37886 37154 37938
rect 38894 37886 38946 37938
rect 40910 37886 40962 37938
rect 4734 37774 4786 37826
rect 8542 37774 8594 37826
rect 9886 37774 9938 37826
rect 21422 37774 21474 37826
rect 26910 37774 26962 37826
rect 29262 37774 29314 37826
rect 32958 37774 33010 37826
rect 37998 37774 38050 37826
rect 38558 37774 38610 37826
rect 38782 37774 38834 37826
rect 41246 37774 41298 37826
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 50558 37606 50610 37658
rect 50662 37606 50714 37658
rect 50766 37606 50818 37658
rect 5854 37438 5906 37490
rect 5966 37438 6018 37490
rect 7534 37438 7586 37490
rect 8878 37438 8930 37490
rect 8990 37438 9042 37490
rect 29374 37438 29426 37490
rect 49310 37438 49362 37490
rect 5294 37326 5346 37378
rect 5518 37326 5570 37378
rect 9550 37326 9602 37378
rect 9662 37326 9714 37378
rect 9886 37326 9938 37378
rect 10446 37326 10498 37378
rect 15934 37326 15986 37378
rect 18510 37326 18562 37378
rect 26798 37326 26850 37378
rect 28030 37326 28082 37378
rect 29486 37326 29538 37378
rect 43262 37326 43314 37378
rect 43822 37326 43874 37378
rect 44046 37326 44098 37378
rect 44158 37326 44210 37378
rect 49086 37326 49138 37378
rect 1822 37214 1874 37266
rect 4846 37214 4898 37266
rect 6078 37214 6130 37266
rect 6526 37214 6578 37266
rect 8318 37214 8370 37266
rect 8766 37214 8818 37266
rect 9998 37214 10050 37266
rect 10222 37214 10274 37266
rect 10670 37214 10722 37266
rect 11006 37214 11058 37266
rect 11790 37214 11842 37266
rect 15262 37214 15314 37266
rect 15822 37214 15874 37266
rect 16494 37214 16546 37266
rect 19070 37214 19122 37266
rect 25566 37214 25618 37266
rect 26238 37214 26290 37266
rect 28478 37214 28530 37266
rect 28926 37214 28978 37266
rect 37550 37214 37602 37266
rect 43150 37214 43202 37266
rect 43710 37214 43762 37266
rect 48638 37214 48690 37266
rect 50430 37214 50482 37266
rect 2494 37102 2546 37154
rect 4622 37102 4674 37154
rect 5070 37102 5122 37154
rect 6974 37102 7026 37154
rect 13918 37102 13970 37154
rect 14366 37102 14418 37154
rect 19406 37102 19458 37154
rect 20078 37102 20130 37154
rect 25342 37102 25394 37154
rect 36430 37102 36482 37154
rect 37102 37102 37154 37154
rect 38222 37102 38274 37154
rect 40350 37102 40402 37154
rect 42702 37102 42754 37154
rect 43486 37102 43538 37154
rect 48190 37102 48242 37154
rect 49198 37102 49250 37154
rect 51102 37102 51154 37154
rect 53230 37102 53282 37154
rect 7198 36990 7250 37042
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 5742 36654 5794 36706
rect 9438 36654 9490 36706
rect 5966 36542 6018 36594
rect 18398 36542 18450 36594
rect 18734 36542 18786 36594
rect 28590 36542 28642 36594
rect 38894 36542 38946 36594
rect 48974 36542 49026 36594
rect 51214 36542 51266 36594
rect 6078 36430 6130 36482
rect 9438 36430 9490 36482
rect 15150 36430 15202 36482
rect 15486 36430 15538 36482
rect 17726 36430 17778 36482
rect 18174 36430 18226 36482
rect 18846 36430 18898 36482
rect 19182 36430 19234 36482
rect 21646 36430 21698 36482
rect 28142 36430 28194 36482
rect 28366 36430 28418 36482
rect 30270 36430 30322 36482
rect 38670 36430 38722 36482
rect 39118 36430 39170 36482
rect 46174 36430 46226 36482
rect 50094 36430 50146 36482
rect 50542 36430 50594 36482
rect 50766 36430 50818 36482
rect 9102 36318 9154 36370
rect 15598 36318 15650 36370
rect 16046 36318 16098 36370
rect 22430 36318 22482 36370
rect 30942 36318 30994 36370
rect 36206 36318 36258 36370
rect 39342 36318 39394 36370
rect 46846 36318 46898 36370
rect 50654 36318 50706 36370
rect 51102 36318 51154 36370
rect 4846 36206 4898 36258
rect 10894 36206 10946 36258
rect 20190 36206 20242 36258
rect 24670 36206 24722 36258
rect 29262 36206 29314 36258
rect 33182 36206 33234 36258
rect 33742 36206 33794 36258
rect 35758 36206 35810 36258
rect 37214 36206 37266 36258
rect 39790 36206 39842 36258
rect 51326 36206 51378 36258
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 50558 36038 50610 36090
rect 50662 36038 50714 36090
rect 50766 36038 50818 36090
rect 4846 35870 4898 35922
rect 7534 35870 7586 35922
rect 21870 35870 21922 35922
rect 22318 35870 22370 35922
rect 22878 35870 22930 35922
rect 38894 35870 38946 35922
rect 46286 35870 46338 35922
rect 5518 35758 5570 35810
rect 8318 35758 8370 35810
rect 8430 35758 8482 35810
rect 22542 35758 22594 35810
rect 36542 35758 36594 35810
rect 38446 35758 38498 35810
rect 44494 35758 44546 35810
rect 46622 35758 46674 35810
rect 49758 35758 49810 35810
rect 5630 35646 5682 35698
rect 7870 35646 7922 35698
rect 8542 35646 8594 35698
rect 16270 35646 16322 35698
rect 22206 35646 22258 35698
rect 22654 35646 22706 35698
rect 23102 35646 23154 35698
rect 23326 35646 23378 35698
rect 33070 35646 33122 35698
rect 36878 35646 36930 35698
rect 37326 35646 37378 35698
rect 37886 35646 37938 35698
rect 38222 35646 38274 35698
rect 45278 35646 45330 35698
rect 45950 35646 46002 35698
rect 46286 35646 46338 35698
rect 49422 35646 49474 35698
rect 50654 35646 50706 35698
rect 15822 35534 15874 35586
rect 16606 35534 16658 35586
rect 23774 35534 23826 35586
rect 33854 35534 33906 35586
rect 35982 35534 36034 35586
rect 41582 35534 41634 35586
rect 42366 35534 42418 35586
rect 49086 35534 49138 35586
rect 5518 35422 5570 35474
rect 8990 35422 9042 35474
rect 53006 35422 53058 35474
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 4622 34974 4674 35026
rect 28366 34974 28418 35026
rect 32174 34974 32226 35026
rect 32734 34974 32786 35026
rect 1822 34862 1874 34914
rect 5518 34862 5570 34914
rect 5854 34862 5906 34914
rect 6190 34862 6242 34914
rect 8766 34862 8818 34914
rect 14366 34862 14418 34914
rect 14814 34862 14866 34914
rect 18510 34862 18562 34914
rect 18846 34862 18898 34914
rect 24558 34862 24610 34914
rect 25342 34862 25394 34914
rect 29262 34862 29314 34914
rect 36206 34862 36258 34914
rect 37886 34862 37938 34914
rect 38334 34862 38386 34914
rect 39118 34862 39170 34914
rect 40014 34862 40066 34914
rect 40574 34862 40626 34914
rect 41582 34862 41634 34914
rect 43934 34862 43986 34914
rect 44830 34862 44882 34914
rect 2494 34750 2546 34802
rect 5070 34750 5122 34802
rect 5742 34750 5794 34802
rect 8990 34750 9042 34802
rect 9550 34750 9602 34802
rect 9886 34750 9938 34802
rect 15038 34750 15090 34802
rect 18958 34750 19010 34802
rect 26126 34750 26178 34802
rect 29934 34750 29986 34802
rect 37326 34750 37378 34802
rect 39342 34750 39394 34802
rect 42590 34750 42642 34802
rect 42702 34750 42754 34802
rect 43822 34750 43874 34802
rect 44942 34750 44994 34802
rect 4958 34638 5010 34690
rect 8094 34638 8146 34690
rect 15486 34638 15538 34690
rect 19406 34638 19458 34690
rect 24222 34638 24274 34690
rect 24670 34638 24722 34690
rect 24894 34638 24946 34690
rect 35758 34638 35810 34690
rect 37102 34638 37154 34690
rect 39454 34638 39506 34690
rect 40910 34638 40962 34690
rect 41246 34638 41298 34690
rect 41918 34638 41970 34690
rect 42366 34638 42418 34690
rect 43598 34638 43650 34690
rect 45166 34638 45218 34690
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 50558 34470 50610 34522
rect 50662 34470 50714 34522
rect 50766 34470 50818 34522
rect 4958 34302 5010 34354
rect 5182 34302 5234 34354
rect 5966 34302 6018 34354
rect 25790 34302 25842 34354
rect 28702 34302 28754 34354
rect 38670 34302 38722 34354
rect 39790 34302 39842 34354
rect 43822 34302 43874 34354
rect 49086 34302 49138 34354
rect 49310 34302 49362 34354
rect 18734 34190 18786 34242
rect 30382 34190 30434 34242
rect 42142 34190 42194 34242
rect 49758 34190 49810 34242
rect 5518 34078 5570 34130
rect 5854 34078 5906 34130
rect 6078 34078 6130 34130
rect 6526 34078 6578 34130
rect 10558 34078 10610 34130
rect 13806 34078 13858 34130
rect 15486 34078 15538 34130
rect 20526 34078 20578 34130
rect 25454 34078 25506 34130
rect 25902 34078 25954 34130
rect 26014 34078 26066 34130
rect 30270 34078 30322 34130
rect 30606 34078 30658 34130
rect 38446 34078 38498 34130
rect 38894 34078 38946 34130
rect 39006 34078 39058 34130
rect 39902 34078 39954 34130
rect 41022 34078 41074 34130
rect 42478 34078 42530 34130
rect 42814 34078 42866 34130
rect 43374 34078 43426 34130
rect 43710 34078 43762 34130
rect 45390 34078 45442 34130
rect 48750 34078 48802 34130
rect 50318 34078 50370 34130
rect 5294 33966 5346 34018
rect 11230 33966 11282 34018
rect 13358 33966 13410 34018
rect 18286 33966 18338 34018
rect 19182 33966 19234 34018
rect 21198 33966 21250 34018
rect 23326 33966 23378 34018
rect 24670 33966 24722 34018
rect 30942 33966 30994 34018
rect 36654 33966 36706 34018
rect 38110 33966 38162 34018
rect 38782 33966 38834 34018
rect 41358 33966 41410 34018
rect 46062 33966 46114 34018
rect 48190 33966 48242 34018
rect 49198 33966 49250 34018
rect 49870 33966 49922 34018
rect 51102 33966 51154 34018
rect 53230 33966 53282 34018
rect 39790 33854 39842 33906
rect 43822 33854 43874 33906
rect 49982 33854 50034 33906
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 9214 33518 9266 33570
rect 29598 33518 29650 33570
rect 30158 33518 30210 33570
rect 33182 33518 33234 33570
rect 9550 33406 9602 33458
rect 11678 33406 11730 33458
rect 16718 33406 16770 33458
rect 21422 33406 21474 33458
rect 31054 33406 31106 33458
rect 41694 33406 41746 33458
rect 45502 33406 45554 33458
rect 48414 33406 48466 33458
rect 50430 33406 50482 33458
rect 5742 33294 5794 33346
rect 5966 33294 6018 33346
rect 6302 33294 6354 33346
rect 10446 33294 10498 33346
rect 10894 33294 10946 33346
rect 14702 33294 14754 33346
rect 15038 33294 15090 33346
rect 17950 33294 18002 33346
rect 18846 33294 18898 33346
rect 19406 33294 19458 33346
rect 19966 33294 20018 33346
rect 20862 33294 20914 33346
rect 21198 33294 21250 33346
rect 23214 33294 23266 33346
rect 25902 33294 25954 33346
rect 29710 33294 29762 33346
rect 29934 33294 29986 33346
rect 30718 33294 30770 33346
rect 33854 33294 33906 33346
rect 45614 33294 45666 33346
rect 45950 33294 46002 33346
rect 49870 33294 49922 33346
rect 50542 33294 50594 33346
rect 5630 33182 5682 33234
rect 10110 33182 10162 33234
rect 10670 33182 10722 33234
rect 11230 33182 11282 33234
rect 15262 33182 15314 33234
rect 19518 33182 19570 33234
rect 20526 33182 20578 33234
rect 21646 33182 21698 33234
rect 21870 33182 21922 33234
rect 23550 33182 23602 33234
rect 25566 33182 25618 33234
rect 33294 33182 33346 33234
rect 33518 33182 33570 33234
rect 33742 33182 33794 33234
rect 34302 33182 34354 33234
rect 45390 33182 45442 33234
rect 6414 33070 6466 33122
rect 6638 33070 6690 33122
rect 7982 33070 8034 33122
rect 8318 33070 8370 33122
rect 8766 33070 8818 33122
rect 9438 33070 9490 33122
rect 10222 33070 10274 33122
rect 10894 33070 10946 33122
rect 20638 33070 20690 33122
rect 23438 33070 23490 33122
rect 24110 33070 24162 33122
rect 25678 33070 25730 33122
rect 26350 33070 26402 33122
rect 29598 33070 29650 33122
rect 30270 33070 30322 33122
rect 30494 33070 30546 33122
rect 31054 33070 31106 33122
rect 31278 33070 31330 33122
rect 32846 33070 32898 33122
rect 33070 33070 33122 33122
rect 40686 33070 40738 33122
rect 50318 33070 50370 33122
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 50558 32902 50610 32954
rect 50662 32902 50714 32954
rect 50766 32902 50818 32954
rect 9886 32734 9938 32786
rect 19070 32734 19122 32786
rect 20862 32734 20914 32786
rect 22766 32734 22818 32786
rect 26238 32734 26290 32786
rect 31166 32734 31218 32786
rect 33406 32734 33458 32786
rect 34078 32734 34130 32786
rect 41246 32734 41298 32786
rect 43374 32734 43426 32786
rect 43598 32734 43650 32786
rect 5294 32622 5346 32674
rect 5630 32622 5682 32674
rect 6078 32622 6130 32674
rect 6190 32622 6242 32674
rect 6414 32622 6466 32674
rect 6638 32622 6690 32674
rect 9550 32622 9602 32674
rect 9662 32622 9714 32674
rect 16158 32622 16210 32674
rect 18958 32622 19010 32674
rect 20414 32622 20466 32674
rect 22990 32622 23042 32674
rect 23102 32622 23154 32674
rect 25678 32622 25730 32674
rect 30382 32622 30434 32674
rect 30942 32622 30994 32674
rect 32398 32622 32450 32674
rect 32622 32622 32674 32674
rect 34302 32622 34354 32674
rect 39678 32622 39730 32674
rect 39902 32622 39954 32674
rect 40462 32622 40514 32674
rect 1822 32510 1874 32562
rect 5854 32510 5906 32562
rect 13694 32510 13746 32562
rect 14254 32510 14306 32562
rect 14366 32510 14418 32562
rect 14814 32510 14866 32562
rect 15038 32510 15090 32562
rect 15262 32510 15314 32562
rect 15486 32510 15538 32562
rect 15598 32510 15650 32562
rect 16046 32510 16098 32562
rect 16382 32510 16434 32562
rect 17838 32510 17890 32562
rect 18398 32510 18450 32562
rect 18510 32510 18562 32562
rect 18846 32510 18898 32562
rect 19854 32510 19906 32562
rect 21198 32510 21250 32562
rect 23550 32510 23602 32562
rect 30494 32510 30546 32562
rect 30830 32510 30882 32562
rect 32286 32510 32338 32562
rect 33742 32510 33794 32562
rect 34526 32510 34578 32562
rect 34750 32510 34802 32562
rect 35310 32510 35362 32562
rect 38782 32510 38834 32562
rect 39230 32510 39282 32562
rect 40910 32510 40962 32562
rect 42926 32510 42978 32562
rect 43150 32510 43202 32562
rect 43598 32510 43650 32562
rect 51102 32510 51154 32562
rect 2494 32398 2546 32450
rect 4622 32398 4674 32450
rect 5406 32398 5458 32450
rect 7086 32398 7138 32450
rect 13022 32398 13074 32450
rect 16830 32398 16882 32450
rect 21646 32398 21698 32450
rect 24670 32398 24722 32450
rect 25566 32398 25618 32450
rect 29934 32398 29986 32450
rect 31502 32398 31554 32450
rect 31950 32398 32002 32450
rect 34414 32398 34466 32450
rect 35982 32398 36034 32450
rect 38110 32398 38162 32450
rect 39454 32398 39506 32450
rect 42590 32398 42642 32450
rect 53006 32398 53058 32450
rect 25454 32286 25506 32338
rect 30382 32286 30434 32338
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 5630 31950 5682 32002
rect 34638 31950 34690 32002
rect 4846 31838 4898 31890
rect 9998 31838 10050 31890
rect 11118 31838 11170 31890
rect 14590 31838 14642 31890
rect 19630 31838 19682 31890
rect 28366 31838 28418 31890
rect 29262 31838 29314 31890
rect 45614 31838 45666 31890
rect 47742 31838 47794 31890
rect 6190 31726 6242 31778
rect 9102 31726 9154 31778
rect 9326 31726 9378 31778
rect 17838 31726 17890 31778
rect 23438 31726 23490 31778
rect 23998 31726 24050 31778
rect 24558 31726 24610 31778
rect 25454 31726 25506 31778
rect 37102 31726 37154 31778
rect 39230 31726 39282 31778
rect 39678 31726 39730 31778
rect 39902 31726 39954 31778
rect 40686 31726 40738 31778
rect 41134 31726 41186 31778
rect 42814 31726 42866 31778
rect 43486 31726 43538 31778
rect 43822 31726 43874 31778
rect 44158 31726 44210 31778
rect 44942 31726 44994 31778
rect 49982 31726 50034 31778
rect 50430 31726 50482 31778
rect 50542 31726 50594 31778
rect 50990 31726 51042 31778
rect 6078 31614 6130 31666
rect 6302 31614 6354 31666
rect 6750 31614 6802 31666
rect 10558 31614 10610 31666
rect 10670 31614 10722 31666
rect 23662 31614 23714 31666
rect 26238 31614 26290 31666
rect 7086 31502 7138 31554
rect 8878 31502 8930 31554
rect 9214 31502 9266 31554
rect 9774 31502 9826 31554
rect 9886 31502 9938 31554
rect 10334 31502 10386 31554
rect 20302 31502 20354 31554
rect 24222 31502 24274 31554
rect 24334 31502 24386 31554
rect 24446 31502 24498 31554
rect 25118 31502 25170 31554
rect 31950 31502 32002 31554
rect 33742 31502 33794 31554
rect 34638 31558 34690 31610
rect 34750 31558 34802 31610
rect 38894 31614 38946 31666
rect 40238 31614 40290 31666
rect 42702 31614 42754 31666
rect 49086 31614 49138 31666
rect 51214 31614 51266 31666
rect 35198 31502 35250 31554
rect 37550 31502 37602 31554
rect 39006 31502 39058 31554
rect 42366 31502 42418 31554
rect 48750 31502 48802 31554
rect 50654 31502 50706 31554
rect 51102 31502 51154 31554
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 50558 31334 50610 31386
rect 50662 31334 50714 31386
rect 50766 31334 50818 31386
rect 6526 31166 6578 31218
rect 7198 31166 7250 31218
rect 7534 31166 7586 31218
rect 33182 31166 33234 31218
rect 35758 31166 35810 31218
rect 36654 31166 36706 31218
rect 38670 31166 38722 31218
rect 38894 31166 38946 31218
rect 39230 31166 39282 31218
rect 42814 31166 42866 31218
rect 43262 31166 43314 31218
rect 43486 31166 43538 31218
rect 43822 31166 43874 31218
rect 44382 31166 44434 31218
rect 48190 31166 48242 31218
rect 49198 31166 49250 31218
rect 49422 31166 49474 31218
rect 6302 31054 6354 31106
rect 10558 31054 10610 31106
rect 18622 31054 18674 31106
rect 26014 31054 26066 31106
rect 37550 31054 37602 31106
rect 37774 31054 37826 31106
rect 43710 31054 43762 31106
rect 44046 31054 44098 31106
rect 44830 31054 44882 31106
rect 45054 31054 45106 31106
rect 51102 31054 51154 31106
rect 6974 30942 7026 30994
rect 9662 30942 9714 30994
rect 9998 30942 10050 30994
rect 10222 30942 10274 30994
rect 11230 30942 11282 30994
rect 15598 30942 15650 30994
rect 16158 30942 16210 30994
rect 17950 30942 18002 30994
rect 24670 30942 24722 30994
rect 25230 30942 25282 30994
rect 25566 30942 25618 30994
rect 25790 30942 25842 30994
rect 29374 30942 29426 30994
rect 36206 30942 36258 30994
rect 36430 30942 36482 30994
rect 36878 30942 36930 30994
rect 37886 30942 37938 30994
rect 37998 30942 38050 30994
rect 38110 30942 38162 30994
rect 38558 30942 38610 30994
rect 39118 30942 39170 30994
rect 43038 30942 43090 30994
rect 44718 30942 44770 30994
rect 47966 30942 48018 30994
rect 48750 30942 48802 30994
rect 50430 30942 50482 30994
rect 6414 30830 6466 30882
rect 9550 30830 9602 30882
rect 10446 30830 10498 30882
rect 12014 30830 12066 30882
rect 14142 30830 14194 30882
rect 16270 30830 16322 30882
rect 16718 30830 16770 30882
rect 18174 30830 18226 30882
rect 25902 30830 25954 30882
rect 26462 30830 26514 30882
rect 30158 30830 30210 30882
rect 32398 30830 32450 30882
rect 35198 30830 35250 30882
rect 36542 30830 36594 30882
rect 48974 30830 49026 30882
rect 49310 30830 49362 30882
rect 53230 30830 53282 30882
rect 39230 30718 39282 30770
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 9438 30382 9490 30434
rect 9550 30382 9602 30434
rect 9886 30382 9938 30434
rect 30830 30382 30882 30434
rect 50206 30382 50258 30434
rect 9774 30270 9826 30322
rect 11118 30270 11170 30322
rect 16270 30270 16322 30322
rect 23886 30270 23938 30322
rect 25118 30270 25170 30322
rect 36990 30270 37042 30322
rect 50430 30270 50482 30322
rect 12798 30158 12850 30210
rect 13806 30158 13858 30210
rect 16382 30158 16434 30210
rect 20526 30158 20578 30210
rect 20862 30158 20914 30210
rect 21198 30158 21250 30210
rect 21534 30158 21586 30210
rect 21870 30158 21922 30210
rect 23998 30158 24050 30210
rect 25566 30158 25618 30210
rect 26238 30158 26290 30210
rect 29374 30158 29426 30210
rect 30942 30158 30994 30210
rect 34638 30158 34690 30210
rect 35086 30158 35138 30210
rect 35534 30158 35586 30210
rect 38222 30158 38274 30210
rect 41358 30158 41410 30210
rect 42590 30158 42642 30210
rect 50542 30158 50594 30210
rect 13470 30046 13522 30098
rect 20638 30046 20690 30098
rect 23326 30046 23378 30098
rect 29710 30046 29762 30098
rect 29822 30046 29874 30098
rect 30046 30046 30098 30098
rect 30270 30046 30322 30098
rect 30494 30046 30546 30098
rect 31278 30046 31330 30098
rect 31838 30046 31890 30098
rect 35310 30046 35362 30098
rect 35870 30046 35922 30098
rect 52222 30046 52274 30098
rect 53230 30046 53282 30098
rect 4958 29934 5010 29986
rect 16270 29934 16322 29986
rect 21422 29934 21474 29986
rect 23550 29934 23602 29986
rect 23774 29934 23826 29986
rect 24558 29934 24610 29986
rect 30718 29934 30770 29986
rect 31166 29934 31218 29986
rect 33630 29934 33682 29986
rect 33966 29934 34018 29986
rect 34302 29934 34354 29986
rect 35758 29934 35810 29986
rect 36430 29934 36482 29986
rect 37550 29934 37602 29986
rect 41134 29934 41186 29986
rect 42030 29934 42082 29986
rect 52894 29934 52946 29986
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 50558 29766 50610 29818
rect 50662 29766 50714 29818
rect 50766 29766 50818 29818
rect 5406 29598 5458 29650
rect 6190 29598 6242 29650
rect 7086 29598 7138 29650
rect 7310 29598 7362 29650
rect 7982 29598 8034 29650
rect 13022 29598 13074 29650
rect 13470 29598 13522 29650
rect 23214 29598 23266 29650
rect 34302 29598 34354 29650
rect 37886 29598 37938 29650
rect 39006 29598 39058 29650
rect 4958 29486 5010 29538
rect 6078 29486 6130 29538
rect 20414 29486 20466 29538
rect 22878 29486 22930 29538
rect 33966 29486 34018 29538
rect 38222 29486 38274 29538
rect 38446 29486 38498 29538
rect 39566 29486 39618 29538
rect 40238 29486 40290 29538
rect 40350 29486 40402 29538
rect 41246 29486 41298 29538
rect 41806 29486 41858 29538
rect 42142 29486 42194 29538
rect 44942 29486 44994 29538
rect 51102 29486 51154 29538
rect 1822 29374 1874 29426
rect 5182 29374 5234 29426
rect 5630 29374 5682 29426
rect 6862 29374 6914 29426
rect 7422 29374 7474 29426
rect 7982 29374 8034 29426
rect 8206 29374 8258 29426
rect 12350 29374 12402 29426
rect 14814 29374 14866 29426
rect 15374 29374 15426 29426
rect 17502 29374 17554 29426
rect 17726 29374 17778 29426
rect 18846 29374 18898 29426
rect 19630 29374 19682 29426
rect 29150 29374 29202 29426
rect 39006 29374 39058 29426
rect 39454 29374 39506 29426
rect 39902 29374 39954 29426
rect 40126 29374 40178 29426
rect 44270 29374 44322 29426
rect 50430 29374 50482 29426
rect 2494 29262 2546 29314
rect 4622 29262 4674 29314
rect 5294 29262 5346 29314
rect 7870 29262 7922 29314
rect 10110 29262 10162 29314
rect 15486 29262 15538 29314
rect 15934 29262 15986 29314
rect 18398 29262 18450 29314
rect 22542 29262 22594 29314
rect 26126 29262 26178 29314
rect 28366 29262 28418 29314
rect 29710 29262 29762 29314
rect 42590 29262 42642 29314
rect 47070 29262 47122 29314
rect 53230 29262 53282 29314
rect 6302 29150 6354 29202
rect 38782 29150 38834 29202
rect 39342 29150 39394 29202
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 2494 28814 2546 28866
rect 2830 28814 2882 28866
rect 5630 28814 5682 28866
rect 5742 28814 5794 28866
rect 5966 28814 6018 28866
rect 10222 28814 10274 28866
rect 11118 28814 11170 28866
rect 11454 28814 11506 28866
rect 19630 28814 19682 28866
rect 25230 28814 25282 28866
rect 25566 28814 25618 28866
rect 29374 28814 29426 28866
rect 38110 28814 38162 28866
rect 40574 28814 40626 28866
rect 41022 28814 41074 28866
rect 42926 28814 42978 28866
rect 19182 28702 19234 28754
rect 21422 28702 21474 28754
rect 25790 28702 25842 28754
rect 26910 28702 26962 28754
rect 27358 28702 27410 28754
rect 35758 28702 35810 28754
rect 39230 28702 39282 28754
rect 40574 28702 40626 28754
rect 41022 28702 41074 28754
rect 43486 28702 43538 28754
rect 46510 28702 46562 28754
rect 50878 28702 50930 28754
rect 3278 28590 3330 28642
rect 4622 28590 4674 28642
rect 6190 28590 6242 28642
rect 7870 28590 7922 28642
rect 9886 28590 9938 28642
rect 11902 28590 11954 28642
rect 16830 28590 16882 28642
rect 17278 28590 17330 28642
rect 17838 28590 17890 28642
rect 20302 28590 20354 28642
rect 20638 28590 20690 28642
rect 24334 28590 24386 28642
rect 24894 28590 24946 28642
rect 26238 28590 26290 28642
rect 29934 28590 29986 28642
rect 30158 28590 30210 28642
rect 30494 28590 30546 28642
rect 36206 28590 36258 28642
rect 37550 28590 37602 28642
rect 37774 28590 37826 28642
rect 39902 28590 39954 28642
rect 41918 28590 41970 28642
rect 42478 28590 42530 28642
rect 42926 28590 42978 28642
rect 44046 28590 44098 28642
rect 44942 28590 44994 28642
rect 46958 28590 47010 28642
rect 47070 28590 47122 28642
rect 48078 28590 48130 28642
rect 2606 28478 2658 28530
rect 11342 28478 11394 28530
rect 17390 28478 17442 28530
rect 19518 28478 19570 28530
rect 19630 28478 19682 28530
rect 20414 28478 20466 28530
rect 30382 28478 30434 28530
rect 31390 28478 31442 28530
rect 41806 28478 41858 28530
rect 45166 28478 45218 28530
rect 47182 28478 47234 28530
rect 48750 28478 48802 28530
rect 4958 28366 5010 28418
rect 8206 28366 8258 28418
rect 10110 28366 10162 28418
rect 26462 28366 26514 28418
rect 29486 28366 29538 28418
rect 29710 28366 29762 28418
rect 30942 28366 30994 28418
rect 31726 28366 31778 28418
rect 39566 28366 39618 28418
rect 47630 28366 47682 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 50558 28198 50610 28250
rect 50662 28198 50714 28250
rect 50766 28198 50818 28250
rect 7310 28030 7362 28082
rect 10446 28030 10498 28082
rect 11566 28030 11618 28082
rect 18846 28030 18898 28082
rect 21870 28030 21922 28082
rect 22206 28030 22258 28082
rect 23998 28030 24050 28082
rect 24222 28030 24274 28082
rect 25342 28030 25394 28082
rect 26910 28030 26962 28082
rect 34078 28030 34130 28082
rect 34750 28030 34802 28082
rect 35646 28030 35698 28082
rect 36430 28030 36482 28082
rect 36542 28030 36594 28082
rect 41358 28030 41410 28082
rect 43374 28030 43426 28082
rect 44942 28030 44994 28082
rect 48302 28030 48354 28082
rect 48862 28030 48914 28082
rect 48974 28030 49026 28082
rect 5630 27918 5682 27970
rect 5742 27918 5794 27970
rect 10782 27918 10834 27970
rect 11006 27918 11058 27970
rect 12686 27918 12738 27970
rect 17502 27918 17554 27970
rect 19966 27918 20018 27970
rect 22990 27918 23042 27970
rect 31838 27918 31890 27970
rect 34302 27918 34354 27970
rect 38782 27918 38834 27970
rect 40238 27918 40290 27970
rect 52894 27918 52946 27970
rect 5406 27806 5458 27858
rect 7422 27806 7474 27858
rect 8990 27806 9042 27858
rect 9662 27806 9714 27858
rect 10110 27806 10162 27858
rect 39790 27862 39842 27914
rect 10334 27806 10386 27858
rect 11566 27806 11618 27858
rect 11902 27806 11954 27858
rect 16158 27806 16210 27858
rect 16718 27806 16770 27858
rect 17390 27806 17442 27858
rect 19406 27806 19458 27858
rect 22542 27806 22594 27858
rect 23438 27806 23490 27858
rect 23774 27806 23826 27858
rect 27246 27806 27298 27858
rect 34750 27806 34802 27858
rect 35758 27806 35810 27858
rect 36094 27806 36146 27858
rect 36318 27806 36370 27858
rect 36766 27806 36818 27858
rect 37662 27806 37714 27858
rect 39006 27806 39058 27858
rect 40014 27806 40066 27858
rect 53230 27806 53282 27858
rect 8878 27694 8930 27746
rect 14814 27694 14866 27746
rect 16830 27694 16882 27746
rect 26238 27694 26290 27746
rect 37214 27694 37266 27746
rect 43710 27694 43762 27746
rect 43934 27694 43986 27746
rect 44494 27694 44546 27746
rect 45502 27694 45554 27746
rect 52670 27694 52722 27746
rect 9550 27582 9602 27634
rect 11230 27582 11282 27634
rect 44158 27582 44210 27634
rect 44494 27582 44546 27634
rect 44942 27582 44994 27634
rect 48750 27582 48802 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 5966 27246 6018 27298
rect 6190 27246 6242 27298
rect 29262 27246 29314 27298
rect 29822 27246 29874 27298
rect 44270 27246 44322 27298
rect 4622 27134 4674 27186
rect 5070 27134 5122 27186
rect 6414 27134 6466 27186
rect 10670 27134 10722 27186
rect 11790 27134 11842 27186
rect 17166 27134 17218 27186
rect 24670 27134 24722 27186
rect 30606 27134 30658 27186
rect 31838 27134 31890 27186
rect 33966 27134 34018 27186
rect 35310 27134 35362 27186
rect 39790 27134 39842 27186
rect 42030 27134 42082 27186
rect 1822 27022 1874 27074
rect 7086 27022 7138 27074
rect 10222 27022 10274 27074
rect 10446 27022 10498 27074
rect 10782 27022 10834 27074
rect 11118 27022 11170 27074
rect 19070 27022 19122 27074
rect 19630 27022 19682 27074
rect 19966 27022 20018 27074
rect 20190 27022 20242 27074
rect 23326 27022 23378 27074
rect 24222 27022 24274 27074
rect 25006 27022 25058 27074
rect 25342 27022 25394 27074
rect 25790 27022 25842 27074
rect 29374 27022 29426 27074
rect 29934 27022 29986 27074
rect 31166 27022 31218 27074
rect 34638 27022 34690 27074
rect 35758 27022 35810 27074
rect 39342 27022 39394 27074
rect 41470 27022 41522 27074
rect 42142 27022 42194 27074
rect 42478 27022 42530 27074
rect 43710 27022 43762 27074
rect 43934 27022 43986 27074
rect 44158 27022 44210 27074
rect 2494 26910 2546 26962
rect 6750 26910 6802 26962
rect 9774 26910 9826 26962
rect 9998 26910 10050 26962
rect 12238 26910 12290 26962
rect 18958 26910 19010 26962
rect 19294 26910 19346 26962
rect 19406 26910 19458 26962
rect 22990 26910 23042 26962
rect 23550 26910 23602 26962
rect 24334 26910 24386 26962
rect 25230 26910 25282 26962
rect 28590 26910 28642 26962
rect 29262 26910 29314 26962
rect 29822 26910 29874 26962
rect 30270 26910 30322 26962
rect 30718 26910 30770 26962
rect 34750 26910 34802 26962
rect 40238 26910 40290 26962
rect 43374 26910 43426 26962
rect 5518 26798 5570 26850
rect 9662 26798 9714 26850
rect 19854 26798 19906 26850
rect 30494 26798 30546 26850
rect 35870 26798 35922 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 50558 26630 50610 26682
rect 50662 26630 50714 26682
rect 50766 26630 50818 26682
rect 21982 26462 22034 26514
rect 25790 26462 25842 26514
rect 29822 26462 29874 26514
rect 30270 26462 30322 26514
rect 30606 26462 30658 26514
rect 34414 26462 34466 26514
rect 34750 26462 34802 26514
rect 35310 26462 35362 26514
rect 35982 26462 36034 26514
rect 36094 26462 36146 26514
rect 41134 26462 41186 26514
rect 42366 26462 42418 26514
rect 5294 26350 5346 26402
rect 5630 26350 5682 26402
rect 7758 26350 7810 26402
rect 8766 26350 8818 26402
rect 19742 26350 19794 26402
rect 29374 26350 29426 26402
rect 30830 26350 30882 26402
rect 30942 26350 30994 26402
rect 31502 26350 31554 26402
rect 38894 26350 38946 26402
rect 41022 26350 41074 26402
rect 43710 26350 43762 26402
rect 5854 26238 5906 26290
rect 6302 26238 6354 26290
rect 8094 26238 8146 26290
rect 8430 26238 8482 26290
rect 19070 26238 19122 26290
rect 28814 26238 28866 26290
rect 29598 26238 29650 26290
rect 35758 26238 35810 26290
rect 36206 26238 36258 26290
rect 36318 26238 36370 26290
rect 38782 26238 38834 26290
rect 43262 26238 43314 26290
rect 45054 26238 45106 26290
rect 49422 26238 49474 26290
rect 49646 26238 49698 26290
rect 49870 26238 49922 26290
rect 50430 26238 50482 26290
rect 5406 26126 5458 26178
rect 28030 26126 28082 26178
rect 29486 26126 29538 26178
rect 42926 26126 42978 26178
rect 45838 26126 45890 26178
rect 47966 26126 48018 26178
rect 49534 26126 49586 26178
rect 51102 26126 51154 26178
rect 53230 26126 53282 26178
rect 38894 26014 38946 26066
rect 41246 26014 41298 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 29710 25678 29762 25730
rect 31390 25678 31442 25730
rect 31726 25678 31778 25730
rect 45726 25678 45778 25730
rect 50990 25678 51042 25730
rect 17054 25566 17106 25618
rect 24222 25566 24274 25618
rect 26350 25566 26402 25618
rect 29262 25566 29314 25618
rect 31726 25566 31778 25618
rect 37102 25566 37154 25618
rect 37998 25566 38050 25618
rect 42030 25566 42082 25618
rect 42590 25566 42642 25618
rect 45502 25566 45554 25618
rect 49758 25566 49810 25618
rect 51102 25566 51154 25618
rect 7646 25454 7698 25506
rect 7982 25454 8034 25506
rect 8542 25454 8594 25506
rect 9438 25454 9490 25506
rect 10558 25454 10610 25506
rect 10782 25454 10834 25506
rect 11006 25454 11058 25506
rect 11118 25454 11170 25506
rect 11566 25454 11618 25506
rect 16270 25454 16322 25506
rect 19182 25454 19234 25506
rect 19854 25454 19906 25506
rect 23886 25454 23938 25506
rect 24558 25454 24610 25506
rect 25566 25454 25618 25506
rect 26238 25454 26290 25506
rect 30830 25454 30882 25506
rect 35422 25454 35474 25506
rect 39006 25454 39058 25506
rect 39790 25454 39842 25506
rect 41134 25454 41186 25506
rect 41582 25454 41634 25506
rect 43038 25454 43090 25506
rect 43150 25454 43202 25506
rect 45838 25454 45890 25506
rect 46062 25454 46114 25506
rect 46286 25454 46338 25506
rect 47742 25454 47794 25506
rect 49870 25454 49922 25506
rect 7198 25342 7250 25394
rect 8094 25342 8146 25394
rect 8206 25342 8258 25394
rect 16606 25342 16658 25394
rect 17614 25342 17666 25394
rect 25230 25342 25282 25394
rect 26014 25342 26066 25394
rect 29822 25342 29874 25394
rect 31166 25342 31218 25394
rect 39342 25342 39394 25394
rect 39678 25342 39730 25394
rect 48190 25342 48242 25394
rect 48414 25342 48466 25394
rect 48750 25342 48802 25394
rect 49086 25342 49138 25394
rect 49310 25342 49362 25394
rect 49646 25342 49698 25394
rect 50206 25342 50258 25394
rect 53230 25342 53282 25394
rect 6078 25230 6130 25282
rect 6414 25230 6466 25282
rect 9886 25230 9938 25282
rect 11118 25230 11170 25282
rect 11902 25230 11954 25282
rect 19518 25230 19570 25282
rect 19742 25230 19794 25282
rect 20302 25230 20354 25282
rect 29710 25230 29762 25282
rect 30382 25230 30434 25282
rect 31054 25230 31106 25282
rect 37550 25230 37602 25282
rect 38558 25230 38610 25282
rect 40014 25230 40066 25282
rect 42254 25230 42306 25282
rect 44046 25230 44098 25282
rect 48078 25230 48130 25282
rect 48862 25230 48914 25282
rect 51214 25230 51266 25282
rect 52894 25230 52946 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 50558 25062 50610 25114
rect 50662 25062 50714 25114
rect 50766 25062 50818 25114
rect 17502 24894 17554 24946
rect 19742 24894 19794 24946
rect 20526 24894 20578 24946
rect 21086 24894 21138 24946
rect 21870 24894 21922 24946
rect 22318 24894 22370 24946
rect 24670 24894 24722 24946
rect 25790 24894 25842 24946
rect 26798 24894 26850 24946
rect 29150 24894 29202 24946
rect 32174 24894 32226 24946
rect 33294 24894 33346 24946
rect 46174 24894 46226 24946
rect 46286 24894 46338 24946
rect 49310 24894 49362 24946
rect 49534 24894 49586 24946
rect 49870 24894 49922 24946
rect 4734 24782 4786 24834
rect 5070 24782 5122 24834
rect 5406 24782 5458 24834
rect 10670 24782 10722 24834
rect 11902 24782 11954 24834
rect 16830 24782 16882 24834
rect 18958 24782 19010 24834
rect 19518 24782 19570 24834
rect 20638 24782 20690 24834
rect 22206 24782 22258 24834
rect 22878 24782 22930 24834
rect 22990 24782 23042 24834
rect 28926 24782 28978 24834
rect 32286 24782 32338 24834
rect 39230 24782 39282 24834
rect 39902 24782 39954 24834
rect 43262 24782 43314 24834
rect 50094 24782 50146 24834
rect 11118 24670 11170 24722
rect 14478 24670 14530 24722
rect 16158 24670 16210 24722
rect 16718 24670 16770 24722
rect 18062 24670 18114 24722
rect 19854 24670 19906 24722
rect 20078 24670 20130 24722
rect 20302 24670 20354 24722
rect 22654 24670 22706 24722
rect 28814 24670 28866 24722
rect 31166 24670 31218 24722
rect 31390 24670 31442 24722
rect 33182 24670 33234 24722
rect 33854 24670 33906 24722
rect 37102 24670 37154 24722
rect 37774 24670 37826 24722
rect 38558 24670 38610 24722
rect 39454 24670 39506 24722
rect 40014 24670 40066 24722
rect 42254 24670 42306 24722
rect 43486 24670 43538 24722
rect 45726 24670 45778 24722
rect 46398 24670 46450 24722
rect 49646 24670 49698 24722
rect 50206 24670 50258 24722
rect 53230 24670 53282 24722
rect 10110 24558 10162 24610
rect 10782 24558 10834 24610
rect 14030 24558 14082 24610
rect 14366 24558 14418 24610
rect 18398 24558 18450 24610
rect 23438 24558 23490 24610
rect 26238 24558 26290 24610
rect 34526 24558 34578 24610
rect 36654 24558 36706 24610
rect 40238 24558 40290 24610
rect 43150 24558 43202 24610
rect 43934 24558 43986 24610
rect 49086 24558 49138 24610
rect 50654 24558 50706 24610
rect 10446 24446 10498 24498
rect 22318 24446 22370 24498
rect 31726 24446 31778 24498
rect 32174 24446 32226 24498
rect 33294 24446 33346 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 34302 24110 34354 24162
rect 45726 24110 45778 24162
rect 4622 23998 4674 24050
rect 5070 23998 5122 24050
rect 6526 23998 6578 24050
rect 7422 23998 7474 24050
rect 8766 23998 8818 24050
rect 17726 23998 17778 24050
rect 19966 23998 20018 24050
rect 24670 23998 24722 24050
rect 26126 23998 26178 24050
rect 28478 23998 28530 24050
rect 40798 23998 40850 24050
rect 47070 23998 47122 24050
rect 1822 23886 1874 23938
rect 5742 23886 5794 23938
rect 7646 23886 7698 23938
rect 8878 23886 8930 23938
rect 15710 23886 15762 23938
rect 20750 23886 20802 23938
rect 21646 23886 21698 23938
rect 25678 23886 25730 23938
rect 31278 23886 31330 23938
rect 31838 23886 31890 23938
rect 34190 23886 34242 23938
rect 37662 23886 37714 23938
rect 39118 23886 39170 23938
rect 41358 23886 41410 23938
rect 43150 23886 43202 23938
rect 46174 23886 46226 23938
rect 2494 23774 2546 23826
rect 5854 23774 5906 23826
rect 6190 23774 6242 23826
rect 6862 23774 6914 23826
rect 8206 23774 8258 23826
rect 8766 23774 8818 23826
rect 9326 23774 9378 23826
rect 15374 23774 15426 23826
rect 22430 23774 22482 23826
rect 27918 23774 27970 23826
rect 28030 23774 28082 23826
rect 33966 23774 34018 23826
rect 34414 23774 34466 23826
rect 34638 23774 34690 23826
rect 34862 23774 34914 23826
rect 34974 23774 35026 23826
rect 37998 23774 38050 23826
rect 38782 23774 38834 23826
rect 38894 23774 38946 23826
rect 42590 23774 42642 23826
rect 43598 23774 43650 23826
rect 44046 23774 44098 23826
rect 45614 23774 45666 23826
rect 5966 23662 6018 23714
rect 6638 23662 6690 23714
rect 7982 23662 8034 23714
rect 8318 23662 8370 23714
rect 9102 23662 9154 23714
rect 25230 23662 25282 23714
rect 26686 23662 26738 23714
rect 27694 23662 27746 23714
rect 30942 23662 30994 23714
rect 32174 23662 32226 23714
rect 32958 23662 33010 23714
rect 37438 23662 37490 23714
rect 37774 23662 37826 23714
rect 43486 23662 43538 23714
rect 45390 23662 45442 23714
rect 45726 23662 45778 23714
rect 46734 23662 46786 23714
rect 47630 23662 47682 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 50558 23494 50610 23546
rect 50662 23494 50714 23546
rect 50766 23494 50818 23546
rect 2606 23326 2658 23378
rect 4734 23326 4786 23378
rect 5406 23326 5458 23378
rect 5630 23326 5682 23378
rect 9774 23326 9826 23378
rect 10558 23326 10610 23378
rect 12350 23326 12402 23378
rect 19294 23326 19346 23378
rect 22542 23326 22594 23378
rect 31166 23326 31218 23378
rect 31502 23326 31554 23378
rect 31838 23326 31890 23378
rect 35198 23326 35250 23378
rect 48862 23326 48914 23378
rect 49086 23326 49138 23378
rect 2830 23214 2882 23266
rect 4510 23214 4562 23266
rect 4958 23214 5010 23266
rect 5854 23214 5906 23266
rect 6190 23214 6242 23266
rect 7646 23214 7698 23266
rect 9550 23214 9602 23266
rect 30830 23214 30882 23266
rect 34750 23214 34802 23266
rect 37662 23214 37714 23266
rect 39342 23214 39394 23266
rect 39566 23214 39618 23266
rect 41694 23214 41746 23266
rect 42030 23214 42082 23266
rect 49758 23214 49810 23266
rect 6302 23102 6354 23154
rect 7198 23102 7250 23154
rect 7870 23102 7922 23154
rect 8430 23102 8482 23154
rect 8654 23102 8706 23154
rect 9998 23102 10050 23154
rect 10222 23102 10274 23154
rect 10782 23102 10834 23154
rect 12686 23102 12738 23154
rect 22318 23102 22370 23154
rect 22654 23102 22706 23154
rect 22990 23102 23042 23154
rect 26462 23102 26514 23154
rect 36654 23102 36706 23154
rect 38110 23102 38162 23154
rect 38446 23102 38498 23154
rect 39230 23102 39282 23154
rect 40014 23102 40066 23154
rect 42814 23102 42866 23154
rect 43038 23102 43090 23154
rect 44158 23102 44210 23154
rect 45726 23102 45778 23154
rect 48750 23102 48802 23154
rect 49310 23102 49362 23154
rect 49870 23102 49922 23154
rect 50430 23102 50482 23154
rect 2494 22990 2546 23042
rect 3278 22990 3330 23042
rect 5742 22990 5794 23042
rect 7422 22990 7474 23042
rect 8990 22990 9042 23042
rect 9886 22990 9938 23042
rect 11342 22990 11394 23042
rect 13470 22990 13522 23042
rect 15598 22990 15650 23042
rect 20974 22990 21026 23042
rect 26126 22990 26178 23042
rect 27246 22990 27298 23042
rect 29374 22990 29426 23042
rect 37214 22990 37266 23042
rect 42142 22990 42194 23042
rect 42702 22990 42754 23042
rect 44494 22990 44546 23042
rect 45278 22990 45330 23042
rect 47966 22990 48018 23042
rect 49534 22990 49586 23042
rect 51102 22990 51154 23042
rect 53230 22990 53282 23042
rect 5070 22878 5122 22930
rect 8878 22878 8930 22930
rect 34750 22878 34802 22930
rect 35198 22878 35250 22930
rect 42590 22878 42642 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 42814 22542 42866 22594
rect 48862 22542 48914 22594
rect 50878 22542 50930 22594
rect 9214 22430 9266 22482
rect 25118 22430 25170 22482
rect 26462 22430 26514 22482
rect 35870 22430 35922 22482
rect 37998 22430 38050 22482
rect 38670 22430 38722 22482
rect 43262 22430 43314 22482
rect 48078 22430 48130 22482
rect 49534 22430 49586 22482
rect 51102 22430 51154 22482
rect 4734 22318 4786 22370
rect 5630 22318 5682 22370
rect 5854 22318 5906 22370
rect 6078 22318 6130 22370
rect 27918 22318 27970 22370
rect 28254 22318 28306 22370
rect 29150 22318 29202 22370
rect 33966 22318 34018 22370
rect 34190 22318 34242 22370
rect 34638 22318 34690 22370
rect 35086 22318 35138 22370
rect 36990 22318 37042 22370
rect 40350 22318 40402 22370
rect 41246 22318 41298 22370
rect 41694 22318 41746 22370
rect 42478 22318 42530 22370
rect 42702 22318 42754 22370
rect 45726 22318 45778 22370
rect 48974 22318 49026 22370
rect 49310 22318 49362 22370
rect 49870 22318 49922 22370
rect 51214 22318 51266 22370
rect 5070 22206 5122 22258
rect 6638 22206 6690 22258
rect 21422 22206 21474 22258
rect 27694 22206 27746 22258
rect 29374 22206 29426 22258
rect 29486 22206 29538 22258
rect 35422 22206 35474 22258
rect 35534 22206 35586 22258
rect 37326 22206 37378 22258
rect 42366 22206 42418 22258
rect 45390 22206 45442 22258
rect 49758 22206 49810 22258
rect 50206 22206 50258 22258
rect 50430 22206 50482 22258
rect 50542 22206 50594 22258
rect 53230 22206 53282 22258
rect 5742 22094 5794 22146
rect 21758 22094 21810 22146
rect 23998 22094 24050 22146
rect 24334 22094 24386 22146
rect 24670 22094 24722 22146
rect 25566 22094 25618 22146
rect 25902 22094 25954 22146
rect 26910 22094 26962 22146
rect 28030 22094 28082 22146
rect 34078 22094 34130 22146
rect 35310 22094 35362 22146
rect 37102 22094 37154 22146
rect 43822 22094 43874 22146
rect 44270 22094 44322 22146
rect 45054 22094 45106 22146
rect 48862 22094 48914 22146
rect 52894 22094 52946 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 50558 21926 50610 21978
rect 50662 21926 50714 21978
rect 50766 21926 50818 21978
rect 5294 21758 5346 21810
rect 5742 21758 5794 21810
rect 8094 21758 8146 21810
rect 8318 21758 8370 21810
rect 9662 21758 9714 21810
rect 13470 21758 13522 21810
rect 14030 21758 14082 21810
rect 21870 21758 21922 21810
rect 22654 21758 22706 21810
rect 34862 21758 34914 21810
rect 38558 21758 38610 21810
rect 41694 21758 41746 21810
rect 43598 21758 43650 21810
rect 46398 21758 46450 21810
rect 49086 21758 49138 21810
rect 49422 21758 49474 21810
rect 49982 21758 50034 21810
rect 53342 21758 53394 21810
rect 2494 21646 2546 21698
rect 23550 21646 23602 21698
rect 23886 21646 23938 21698
rect 33854 21646 33906 21698
rect 35982 21646 36034 21698
rect 40014 21646 40066 21698
rect 44046 21646 44098 21698
rect 47966 21646 48018 21698
rect 48750 21646 48802 21698
rect 48862 21646 48914 21698
rect 49310 21646 49362 21698
rect 1822 21534 1874 21586
rect 7982 21534 8034 21586
rect 10446 21534 10498 21586
rect 19630 21534 19682 21586
rect 20078 21534 20130 21586
rect 20638 21534 20690 21586
rect 21534 21534 21586 21586
rect 23214 21534 23266 21586
rect 33182 21534 33234 21586
rect 33518 21534 33570 21586
rect 35310 21534 35362 21586
rect 40238 21534 40290 21586
rect 40910 21534 40962 21586
rect 41134 21534 41186 21586
rect 43934 21534 43986 21586
rect 45838 21534 45890 21586
rect 47294 21534 47346 21586
rect 47630 21534 47682 21586
rect 49646 21534 49698 21586
rect 4622 21422 4674 21474
rect 8654 21422 8706 21474
rect 9998 21422 10050 21474
rect 11230 21422 11282 21474
rect 15038 21422 15090 21474
rect 15598 21422 15650 21474
rect 19182 21422 19234 21474
rect 22318 21422 22370 21474
rect 33406 21422 33458 21474
rect 38110 21422 38162 21474
rect 39566 21422 39618 21474
rect 42142 21422 42194 21474
rect 44494 21422 44546 21474
rect 44942 21422 44994 21474
rect 45390 21422 45442 21474
rect 46734 21422 46786 21474
rect 50430 21422 50482 21474
rect 10110 21310 10162 21362
rect 41246 21310 41298 21362
rect 44270 21310 44322 21362
rect 44942 21310 44994 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 7534 20974 7586 21026
rect 10446 20974 10498 21026
rect 42814 20974 42866 21026
rect 14590 20862 14642 20914
rect 18510 20862 18562 20914
rect 20414 20862 20466 20914
rect 29822 20862 29874 20914
rect 31726 20862 31778 20914
rect 33854 20862 33906 20914
rect 39230 20862 39282 20914
rect 41022 20862 41074 20914
rect 43486 20862 43538 20914
rect 45390 20862 45442 20914
rect 49982 20862 50034 20914
rect 9998 20750 10050 20802
rect 10222 20750 10274 20802
rect 10558 20750 10610 20802
rect 14142 20750 14194 20802
rect 14814 20750 14866 20802
rect 15598 20750 15650 20802
rect 19070 20750 19122 20802
rect 19966 20750 20018 20802
rect 22206 20750 22258 20802
rect 27022 20750 27074 20802
rect 27694 20750 27746 20802
rect 27918 20750 27970 20802
rect 28254 20750 28306 20802
rect 28478 20750 28530 20802
rect 29374 20750 29426 20802
rect 30270 20750 30322 20802
rect 30606 20750 30658 20802
rect 30942 20750 30994 20802
rect 41582 20750 41634 20802
rect 43038 20750 43090 20802
rect 43262 20750 43314 20802
rect 45950 20750 46002 20802
rect 46510 20750 46562 20802
rect 7870 20638 7922 20690
rect 13806 20638 13858 20690
rect 14478 20638 14530 20690
rect 15262 20638 15314 20690
rect 16382 20638 16434 20690
rect 18846 20638 18898 20690
rect 19630 20638 19682 20690
rect 27246 20638 27298 20690
rect 29038 20638 29090 20690
rect 43822 20638 43874 20690
rect 44942 20638 44994 20690
rect 7646 20526 7698 20578
rect 10782 20526 10834 20578
rect 21870 20526 21922 20578
rect 27358 20526 27410 20578
rect 28366 20526 28418 20578
rect 29262 20526 29314 20578
rect 30494 20526 30546 20578
rect 42366 20526 42418 20578
rect 44158 20526 44210 20578
rect 44830 20526 44882 20578
rect 46958 20526 47010 20578
rect 47406 20526 47458 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 50558 20358 50610 20410
rect 50662 20358 50714 20410
rect 50766 20358 50818 20410
rect 9886 20190 9938 20242
rect 18846 20190 18898 20242
rect 28366 20190 28418 20242
rect 28478 20190 28530 20242
rect 30046 20190 30098 20242
rect 6862 20078 6914 20130
rect 8654 20078 8706 20130
rect 15150 20078 15202 20130
rect 15822 20078 15874 20130
rect 18510 20078 18562 20130
rect 24782 20078 24834 20130
rect 25790 20078 25842 20130
rect 28142 20078 28194 20130
rect 28702 20078 28754 20130
rect 30606 20078 30658 20130
rect 42702 20078 42754 20130
rect 44718 20078 44770 20130
rect 49758 20078 49810 20130
rect 6414 19966 6466 20018
rect 7086 19966 7138 20018
rect 7310 19966 7362 20018
rect 8318 19966 8370 20018
rect 8990 19966 9042 20018
rect 10110 19966 10162 20018
rect 14926 19966 14978 20018
rect 15486 19966 15538 20018
rect 16158 19966 16210 20018
rect 25230 19966 25282 20018
rect 25566 19966 25618 20018
rect 28030 19966 28082 20018
rect 28814 19966 28866 20018
rect 40126 19966 40178 20018
rect 40350 19966 40402 20018
rect 41358 19966 41410 20018
rect 43710 19966 43762 20018
rect 44158 19966 44210 20018
rect 46286 19966 46338 20018
rect 49198 19966 49250 20018
rect 49534 19966 49586 20018
rect 50430 19966 50482 20018
rect 8094 19854 8146 19906
rect 9774 19854 9826 19906
rect 16606 19854 16658 19906
rect 25342 19854 25394 19906
rect 27694 19854 27746 19906
rect 29262 19854 29314 19906
rect 40910 19854 40962 19906
rect 45502 19854 45554 19906
rect 46846 19854 46898 19906
rect 49646 19854 49698 19906
rect 51102 19854 51154 19906
rect 53230 19854 53282 19906
rect 7982 19742 8034 19794
rect 39790 19742 39842 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 4958 19406 5010 19458
rect 7086 19406 7138 19458
rect 11454 19406 11506 19458
rect 38446 19406 38498 19458
rect 51102 19406 51154 19458
rect 8542 19294 8594 19346
rect 11230 19294 11282 19346
rect 12014 19294 12066 19346
rect 15374 19294 15426 19346
rect 18622 19294 18674 19346
rect 23998 19294 24050 19346
rect 26126 19294 26178 19346
rect 30830 19294 30882 19346
rect 31166 19294 31218 19346
rect 39454 19294 39506 19346
rect 41694 19294 41746 19346
rect 45950 19294 46002 19346
rect 5630 19182 5682 19234
rect 5854 19182 5906 19234
rect 7086 19182 7138 19234
rect 7982 19182 8034 19234
rect 8990 19182 9042 19234
rect 11006 19182 11058 19234
rect 15710 19182 15762 19234
rect 23214 19182 23266 19234
rect 30494 19182 30546 19234
rect 31502 19182 31554 19234
rect 32174 19182 32226 19234
rect 32510 19182 32562 19234
rect 33294 19182 33346 19234
rect 34302 19182 34354 19234
rect 34862 19182 34914 19234
rect 39790 19182 39842 19234
rect 46286 19182 46338 19234
rect 47966 19182 48018 19234
rect 49534 19182 49586 19234
rect 49758 19182 49810 19234
rect 49982 19182 50034 19234
rect 53230 19182 53282 19234
rect 5070 19070 5122 19122
rect 6526 19070 6578 19122
rect 6750 19070 6802 19122
rect 7646 19070 7698 19122
rect 10110 19070 10162 19122
rect 11566 19070 11618 19122
rect 16494 19070 16546 19122
rect 22766 19070 22818 19122
rect 22878 19070 22930 19122
rect 31614 19070 31666 19122
rect 31838 19070 31890 19122
rect 32846 19070 32898 19122
rect 34638 19070 34690 19122
rect 35198 19070 35250 19122
rect 35310 19070 35362 19122
rect 38670 19070 38722 19122
rect 39118 19070 39170 19122
rect 46622 19070 46674 19122
rect 48526 19070 48578 19122
rect 48862 19070 48914 19122
rect 49198 19070 49250 19122
rect 50206 19070 50258 19122
rect 50318 19070 50370 19122
rect 50766 19070 50818 19122
rect 50990 19070 51042 19122
rect 52894 19070 52946 19122
rect 4958 18958 5010 19010
rect 6190 18958 6242 19010
rect 6638 18958 6690 19010
rect 10446 18958 10498 19010
rect 22318 18958 22370 19010
rect 22542 18958 22594 19010
rect 32622 18958 32674 19010
rect 32734 18958 32786 19010
rect 33966 18958 34018 19010
rect 34414 18958 34466 19010
rect 34974 18958 35026 19010
rect 35086 18958 35138 19010
rect 38558 18958 38610 19010
rect 42142 18958 42194 19010
rect 48190 18958 48242 19010
rect 49310 18958 49362 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 50558 18790 50610 18842
rect 50662 18790 50714 18842
rect 50766 18790 50818 18842
rect 7646 18622 7698 18674
rect 15150 18622 15202 18674
rect 25118 18622 25170 18674
rect 29262 18622 29314 18674
rect 38334 18622 38386 18674
rect 51102 18622 51154 18674
rect 53342 18622 53394 18674
rect 6414 18510 6466 18562
rect 18510 18510 18562 18562
rect 25342 18510 25394 18562
rect 45502 18510 45554 18562
rect 45838 18510 45890 18562
rect 50094 18510 50146 18562
rect 1822 18398 1874 18450
rect 2494 18398 2546 18450
rect 5518 18398 5570 18450
rect 5966 18398 6018 18450
rect 6302 18398 6354 18450
rect 6638 18398 6690 18450
rect 11902 18398 11954 18450
rect 19854 18398 19906 18450
rect 25454 18398 25506 18450
rect 26238 18398 26290 18450
rect 27022 18398 27074 18450
rect 35422 18398 35474 18450
rect 36094 18398 36146 18450
rect 38894 18398 38946 18450
rect 41806 18398 41858 18450
rect 42254 18398 42306 18450
rect 46734 18398 46786 18450
rect 49870 18398 49922 18450
rect 50542 18398 50594 18450
rect 4622 18286 4674 18338
rect 5070 18286 5122 18338
rect 12574 18286 12626 18338
rect 14702 18286 14754 18338
rect 20638 18286 20690 18338
rect 22766 18286 22818 18338
rect 23214 18286 23266 18338
rect 25902 18286 25954 18338
rect 33182 18286 33234 18338
rect 42926 18286 42978 18338
rect 45054 18286 45106 18338
rect 46174 18286 46226 18338
rect 47182 18286 47234 18338
rect 50318 18286 50370 18338
rect 50878 18286 50930 18338
rect 51102 18286 51154 18338
rect 18398 18174 18450 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 34078 17838 34130 17890
rect 6526 17726 6578 17778
rect 15710 17726 15762 17778
rect 21422 17726 21474 17778
rect 30718 17726 30770 17778
rect 36430 17726 36482 17778
rect 49422 17726 49474 17778
rect 6750 17614 6802 17666
rect 21870 17614 21922 17666
rect 29598 17614 29650 17666
rect 30046 17614 30098 17666
rect 33966 17614 34018 17666
rect 37662 17614 37714 17666
rect 37998 17614 38050 17666
rect 38110 17614 38162 17666
rect 39118 17614 39170 17666
rect 40462 17614 40514 17666
rect 42254 17614 42306 17666
rect 43262 17614 43314 17666
rect 48526 17614 48578 17666
rect 49310 17614 49362 17666
rect 49870 17614 49922 17666
rect 6302 17502 6354 17554
rect 6414 17502 6466 17554
rect 6526 17502 6578 17554
rect 7982 17502 8034 17554
rect 15150 17502 15202 17554
rect 21310 17502 21362 17554
rect 21646 17502 21698 17554
rect 23550 17502 23602 17554
rect 23662 17502 23714 17554
rect 33406 17502 33458 17554
rect 38558 17502 38610 17554
rect 42030 17502 42082 17554
rect 47630 17502 47682 17554
rect 48190 17502 48242 17554
rect 48302 17502 48354 17554
rect 49646 17502 49698 17554
rect 4846 17390 4898 17442
rect 7646 17390 7698 17442
rect 15262 17390 15314 17442
rect 23326 17390 23378 17442
rect 32958 17390 33010 17442
rect 33518 17390 33570 17442
rect 36318 17390 36370 17442
rect 40014 17390 40066 17442
rect 42926 17390 42978 17442
rect 47742 17390 47794 17442
rect 47966 17390 48018 17442
rect 48862 17390 48914 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 50558 17222 50610 17274
rect 50662 17222 50714 17274
rect 50766 17222 50818 17274
rect 4622 17054 4674 17106
rect 12910 17054 12962 17106
rect 16606 17054 16658 17106
rect 18174 17054 18226 17106
rect 34526 17054 34578 17106
rect 34750 17054 34802 17106
rect 36318 17054 36370 17106
rect 36542 17054 36594 17106
rect 38110 17054 38162 17106
rect 38334 17054 38386 17106
rect 39006 17054 39058 17106
rect 41246 17054 41298 17106
rect 41918 17054 41970 17106
rect 50094 17054 50146 17106
rect 4734 16942 4786 16994
rect 13022 16942 13074 16994
rect 14478 16942 14530 16994
rect 16046 16942 16098 16994
rect 19294 16942 19346 16994
rect 33742 16942 33794 16994
rect 35422 16942 35474 16994
rect 37102 16942 37154 16994
rect 42702 16942 42754 16994
rect 42814 16942 42866 16994
rect 48862 16942 48914 16994
rect 49758 16942 49810 16994
rect 49870 16942 49922 16994
rect 51102 16942 51154 16994
rect 9662 16830 9714 16882
rect 12798 16830 12850 16882
rect 13246 16830 13298 16882
rect 13470 16830 13522 16882
rect 14590 16830 14642 16882
rect 14814 16830 14866 16882
rect 15262 16830 15314 16882
rect 15822 16830 15874 16882
rect 16606 16830 16658 16882
rect 17390 16830 17442 16882
rect 17726 16830 17778 16882
rect 18174 16830 18226 16882
rect 18622 16830 18674 16882
rect 24110 16830 24162 16882
rect 33406 16830 33458 16882
rect 34302 16830 34354 16882
rect 35310 16830 35362 16882
rect 36430 16830 36482 16882
rect 37550 16830 37602 16882
rect 37886 16830 37938 16882
rect 41582 16830 41634 16882
rect 42030 16830 42082 16882
rect 42366 16830 42418 16882
rect 48750 16830 48802 16882
rect 49086 16830 49138 16882
rect 49422 16830 49474 16882
rect 50318 16830 50370 16882
rect 10334 16718 10386 16770
rect 12462 16718 12514 16770
rect 21422 16718 21474 16770
rect 22318 16718 22370 16770
rect 25342 16718 25394 16770
rect 53230 16718 53282 16770
rect 4510 16606 4562 16658
rect 15038 16606 15090 16658
rect 16382 16606 16434 16658
rect 17838 16606 17890 16658
rect 25118 16606 25170 16658
rect 25342 16606 25394 16658
rect 41806 16606 41858 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 6414 16270 6466 16322
rect 10446 16270 10498 16322
rect 11678 16270 11730 16322
rect 15262 16270 15314 16322
rect 16494 16270 16546 16322
rect 32958 16270 33010 16322
rect 4622 16158 4674 16210
rect 5070 16158 5122 16210
rect 18174 16158 18226 16210
rect 21646 16158 21698 16210
rect 25566 16158 25618 16210
rect 26014 16158 26066 16210
rect 40462 16158 40514 16210
rect 44830 16158 44882 16210
rect 1822 16046 1874 16098
rect 5966 16046 6018 16098
rect 6190 16046 6242 16098
rect 7310 16046 7362 16098
rect 7534 16046 7586 16098
rect 7982 16046 8034 16098
rect 9886 16046 9938 16098
rect 10110 16046 10162 16098
rect 10558 16046 10610 16098
rect 11790 16046 11842 16098
rect 16270 16046 16322 16098
rect 16718 16046 16770 16098
rect 17502 16046 17554 16098
rect 17726 16046 17778 16098
rect 22654 16046 22706 16098
rect 32846 16046 32898 16098
rect 37998 16046 38050 16098
rect 38558 16046 38610 16098
rect 38670 16046 38722 16098
rect 40014 16046 40066 16098
rect 40798 16046 40850 16098
rect 42590 16046 42642 16098
rect 47742 16046 47794 16098
rect 48190 16046 48242 16098
rect 48862 16046 48914 16098
rect 49646 16046 49698 16098
rect 50206 16046 50258 16098
rect 53118 16046 53170 16098
rect 2494 15934 2546 15986
rect 6526 15934 6578 15986
rect 15374 15934 15426 15986
rect 15598 15934 15650 15986
rect 16942 15934 16994 15986
rect 17390 15934 17442 15986
rect 23438 15934 23490 15986
rect 34862 15934 34914 15986
rect 38334 15934 38386 15986
rect 39678 15934 39730 15986
rect 40686 15934 40738 15986
rect 42926 15934 42978 15986
rect 46958 15934 47010 15986
rect 48638 15934 48690 15986
rect 49870 15934 49922 15986
rect 52894 15934 52946 15986
rect 7422 15822 7474 15874
rect 10222 15822 10274 15874
rect 12686 15822 12738 15874
rect 16494 15822 16546 15874
rect 37102 15822 37154 15874
rect 37774 15822 37826 15874
rect 42814 15822 42866 15874
rect 48526 15822 48578 15874
rect 50094 15822 50146 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 50558 15654 50610 15706
rect 50662 15654 50714 15706
rect 50766 15654 50818 15706
rect 2270 15486 2322 15538
rect 4622 15486 4674 15538
rect 8542 15486 8594 15538
rect 9662 15486 9714 15538
rect 12126 15486 12178 15538
rect 12798 15486 12850 15538
rect 18510 15486 18562 15538
rect 25342 15486 25394 15538
rect 29822 15486 29874 15538
rect 31390 15486 31442 15538
rect 32398 15486 32450 15538
rect 41022 15486 41074 15538
rect 43262 15486 43314 15538
rect 43486 15486 43538 15538
rect 44494 15486 44546 15538
rect 46398 15486 46450 15538
rect 46734 15486 46786 15538
rect 47966 15486 48018 15538
rect 48638 15486 48690 15538
rect 49870 15486 49922 15538
rect 50430 15486 50482 15538
rect 53342 15486 53394 15538
rect 4958 15374 5010 15426
rect 7086 15374 7138 15426
rect 7198 15374 7250 15426
rect 8206 15374 8258 15426
rect 8766 15374 8818 15426
rect 8878 15374 8930 15426
rect 13134 15374 13186 15426
rect 18622 15374 18674 15426
rect 19742 15374 19794 15426
rect 20750 15374 20802 15426
rect 27582 15374 27634 15426
rect 30942 15374 30994 15426
rect 39790 15374 39842 15426
rect 41470 15374 41522 15426
rect 42366 15374 42418 15426
rect 44606 15374 44658 15426
rect 47070 15374 47122 15426
rect 48862 15374 48914 15426
rect 48974 15374 49026 15426
rect 49534 15374 49586 15426
rect 49646 15374 49698 15426
rect 50094 15374 50146 15426
rect 2606 15262 2658 15314
rect 7534 15262 7586 15314
rect 7982 15262 8034 15314
rect 8094 15262 8146 15314
rect 12350 15262 12402 15314
rect 14030 15262 14082 15314
rect 18398 15262 18450 15314
rect 19070 15262 19122 15314
rect 24110 15262 24162 15314
rect 26798 15262 26850 15314
rect 30718 15262 30770 15314
rect 31614 15262 31666 15314
rect 31838 15262 31890 15314
rect 34414 15262 34466 15314
rect 36206 15262 36258 15314
rect 36542 15262 36594 15314
rect 36990 15262 37042 15314
rect 37998 15262 38050 15314
rect 41246 15262 41298 15314
rect 42142 15262 42194 15314
rect 42254 15262 42306 15314
rect 42478 15262 42530 15314
rect 42590 15262 42642 15314
rect 43710 15262 43762 15314
rect 44046 15262 44098 15314
rect 50318 15262 50370 15314
rect 50654 15262 50706 15314
rect 15150 15150 15202 15202
rect 16494 15150 16546 15202
rect 18846 15150 18898 15202
rect 22654 15150 22706 15202
rect 26462 15150 26514 15202
rect 31726 15150 31778 15202
rect 33966 15150 34018 15202
rect 34638 15150 34690 15202
rect 38446 15150 38498 15202
rect 43598 15150 43650 15202
rect 44382 15150 44434 15202
rect 7086 15038 7138 15090
rect 20638 15038 20690 15090
rect 38894 15038 38946 15090
rect 39902 15038 39954 15090
rect 40910 15038 40962 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 19070 14702 19122 14754
rect 31502 14702 31554 14754
rect 33070 14702 33122 14754
rect 35646 14702 35698 14754
rect 15038 14590 15090 14642
rect 23326 14590 23378 14642
rect 34750 14590 34802 14642
rect 41134 14590 41186 14642
rect 52670 14590 52722 14642
rect 6974 14478 7026 14530
rect 7534 14478 7586 14530
rect 10446 14478 10498 14530
rect 11342 14478 11394 14530
rect 12014 14478 12066 14530
rect 16270 14478 16322 14530
rect 16606 14478 16658 14530
rect 17278 14478 17330 14530
rect 19070 14478 19122 14530
rect 22878 14478 22930 14530
rect 25342 14478 25394 14530
rect 31950 14478 32002 14530
rect 32174 14478 32226 14530
rect 32510 14478 32562 14530
rect 35870 14478 35922 14530
rect 38670 14478 38722 14530
rect 38894 14478 38946 14530
rect 40686 14478 40738 14530
rect 41022 14478 41074 14530
rect 41246 14478 41298 14530
rect 43374 14478 43426 14530
rect 46398 14478 46450 14530
rect 48526 14478 48578 14530
rect 48862 14478 48914 14530
rect 49086 14478 49138 14530
rect 11006 14366 11058 14418
rect 18734 14366 18786 14418
rect 23102 14366 23154 14418
rect 23438 14366 23490 14418
rect 25790 14366 25842 14418
rect 31278 14366 31330 14418
rect 32286 14366 32338 14418
rect 33182 14366 33234 14418
rect 35310 14366 35362 14418
rect 39118 14366 39170 14418
rect 41918 14366 41970 14418
rect 43038 14366 43090 14418
rect 46062 14366 46114 14418
rect 7086 14254 7138 14306
rect 7198 14254 7250 14306
rect 8542 14254 8594 14306
rect 10222 14254 10274 14306
rect 11678 14254 11730 14306
rect 16942 14254 16994 14306
rect 17614 14254 17666 14306
rect 25118 14254 25170 14306
rect 26126 14254 26178 14306
rect 26574 14254 26626 14306
rect 31390 14254 31442 14306
rect 32398 14254 32450 14306
rect 33070 14254 33122 14306
rect 40798 14254 40850 14306
rect 42254 14254 42306 14306
rect 46174 14254 46226 14306
rect 46846 14254 46898 14306
rect 48862 14254 48914 14306
rect 52222 14254 52274 14306
rect 53230 14254 53282 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 50558 14086 50610 14138
rect 50662 14086 50714 14138
rect 50766 14086 50818 14138
rect 7310 13918 7362 13970
rect 9550 13918 9602 13970
rect 10334 13918 10386 13970
rect 12574 13918 12626 13970
rect 15598 13918 15650 13970
rect 16942 13918 16994 13970
rect 18622 13918 18674 13970
rect 32286 13918 32338 13970
rect 33854 13918 33906 13970
rect 39678 13918 39730 13970
rect 40014 13918 40066 13970
rect 16158 13806 16210 13858
rect 16382 13806 16434 13858
rect 18286 13806 18338 13858
rect 19630 13806 19682 13858
rect 27918 13806 27970 13858
rect 31838 13806 31890 13858
rect 32510 13806 32562 13858
rect 33630 13806 33682 13858
rect 5182 13694 5234 13746
rect 5966 13694 6018 13746
rect 6190 13694 6242 13746
rect 6414 13694 6466 13746
rect 6638 13694 6690 13746
rect 6974 13694 7026 13746
rect 9774 13694 9826 13746
rect 12350 13694 12402 13746
rect 15822 13694 15874 13746
rect 15934 13694 15986 13746
rect 18510 13694 18562 13746
rect 19070 13694 19122 13746
rect 20302 13694 20354 13746
rect 21534 13694 21586 13746
rect 27134 13694 27186 13746
rect 32062 13694 32114 13746
rect 35534 13694 35586 13746
rect 50318 13694 50370 13746
rect 5070 13582 5122 13634
rect 6078 13582 6130 13634
rect 17614 13582 17666 13634
rect 18734 13582 18786 13634
rect 19518 13582 19570 13634
rect 22206 13582 22258 13634
rect 24334 13582 24386 13634
rect 25342 13582 25394 13634
rect 26798 13582 26850 13634
rect 30046 13582 30098 13634
rect 35758 13582 35810 13634
rect 36206 13582 36258 13634
rect 49982 13582 50034 13634
rect 51102 13582 51154 13634
rect 53230 13582 53282 13634
rect 4846 13470 4898 13522
rect 7086 13470 7138 13522
rect 7422 13470 7474 13522
rect 19406 13470 19458 13522
rect 31950 13470 32002 13522
rect 33966 13470 34018 13522
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 6190 13134 6242 13186
rect 6414 13134 6466 13186
rect 6862 13134 6914 13186
rect 10670 13134 10722 13186
rect 14366 13134 14418 13186
rect 15486 13134 15538 13186
rect 15822 13134 15874 13186
rect 18622 13134 18674 13186
rect 41918 13134 41970 13186
rect 50542 13134 50594 13186
rect 50878 13134 50930 13186
rect 2494 13022 2546 13074
rect 4622 13022 4674 13074
rect 4958 13022 5010 13074
rect 7198 13022 7250 13074
rect 11566 13022 11618 13074
rect 11902 13022 11954 13074
rect 22206 13022 22258 13074
rect 24782 13022 24834 13074
rect 28590 13022 28642 13074
rect 46846 13022 46898 13074
rect 1822 12910 1874 12962
rect 5070 12910 5122 12962
rect 5742 12910 5794 12962
rect 6862 12910 6914 12962
rect 11006 12910 11058 12962
rect 13918 12910 13970 12962
rect 14254 12910 14306 12962
rect 14478 12910 14530 12962
rect 15150 12910 15202 12962
rect 15822 12910 15874 12962
rect 18062 12910 18114 12962
rect 18398 12910 18450 12962
rect 18846 12910 18898 12962
rect 21870 12910 21922 12962
rect 22094 12910 22146 12962
rect 22430 12910 22482 12962
rect 25678 12910 25730 12962
rect 35646 12910 35698 12962
rect 36206 12910 36258 12962
rect 38110 12910 38162 12962
rect 38334 12910 38386 12962
rect 38782 12910 38834 12962
rect 42254 12910 42306 12962
rect 43934 12910 43986 12962
rect 49758 12910 49810 12962
rect 5630 12798 5682 12850
rect 23998 12798 24050 12850
rect 24222 12798 24274 12850
rect 24334 12798 24386 12850
rect 26462 12798 26514 12850
rect 43710 12798 43762 12850
rect 48974 12798 49026 12850
rect 6526 12686 6578 12738
rect 10782 12686 10834 12738
rect 14702 12686 14754 12738
rect 18174 12686 18226 12738
rect 25342 12686 25394 12738
rect 35870 12686 35922 12738
rect 35982 12686 36034 12738
rect 36094 12686 36146 12738
rect 38446 12686 38498 12738
rect 38558 12686 38610 12738
rect 42030 12686 42082 12738
rect 45614 12686 45666 12738
rect 45950 12686 46002 12738
rect 46286 12686 46338 12738
rect 50206 12686 50258 12738
rect 50766 12686 50818 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 50558 12518 50610 12570
rect 50662 12518 50714 12570
rect 50766 12518 50818 12570
rect 10670 12350 10722 12402
rect 14030 12350 14082 12402
rect 24110 12350 24162 12402
rect 27022 12350 27074 12402
rect 27694 12350 27746 12402
rect 28814 12350 28866 12402
rect 41022 12350 41074 12402
rect 45390 12350 45442 12402
rect 45726 12350 45778 12402
rect 48862 12350 48914 12402
rect 9886 12238 9938 12290
rect 12126 12238 12178 12290
rect 13918 12238 13970 12290
rect 14142 12238 14194 12290
rect 14590 12238 14642 12290
rect 14814 12238 14866 12290
rect 27582 12238 27634 12290
rect 36318 12238 36370 12290
rect 36542 12238 36594 12290
rect 48750 12238 48802 12290
rect 48974 12238 49026 12290
rect 52446 12238 52498 12290
rect 8094 12126 8146 12178
rect 10110 12126 10162 12178
rect 10670 12126 10722 12178
rect 12462 12126 12514 12178
rect 12910 12126 12962 12178
rect 13470 12126 13522 12178
rect 21758 12126 21810 12178
rect 21870 12126 21922 12178
rect 22318 12126 22370 12178
rect 23886 12126 23938 12178
rect 24222 12126 24274 12178
rect 26686 12126 26738 12178
rect 26910 12126 26962 12178
rect 27358 12126 27410 12178
rect 29262 12126 29314 12178
rect 35982 12126 36034 12178
rect 37102 12126 37154 12178
rect 41582 12126 41634 12178
rect 4846 12014 4898 12066
rect 7870 12014 7922 12066
rect 12238 12014 12290 12066
rect 14478 12014 14530 12066
rect 19294 12014 19346 12066
rect 22094 12014 22146 12066
rect 24670 12014 24722 12066
rect 29934 12014 29986 12066
rect 32062 12014 32114 12066
rect 33070 12014 33122 12066
rect 35198 12014 35250 12066
rect 36430 12014 36482 12066
rect 37886 12014 37938 12066
rect 40014 12014 40066 12066
rect 42366 12014 42418 12066
rect 44494 12014 44546 12066
rect 46174 12014 46226 12066
rect 52782 12014 52834 12066
rect 53342 12014 53394 12066
rect 8318 11902 8370 11954
rect 8766 11902 8818 11954
rect 10334 11902 10386 11954
rect 12574 11902 12626 11954
rect 19182 11902 19234 11954
rect 27694 11902 27746 11954
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 15598 11566 15650 11618
rect 38110 11566 38162 11618
rect 38446 11566 38498 11618
rect 40462 11566 40514 11618
rect 41022 11566 41074 11618
rect 42030 11566 42082 11618
rect 5854 11454 5906 11506
rect 7870 11454 7922 11506
rect 14478 11454 14530 11506
rect 17726 11454 17778 11506
rect 19854 11454 19906 11506
rect 22206 11454 22258 11506
rect 24334 11454 24386 11506
rect 31838 11454 31890 11506
rect 41246 11454 41298 11506
rect 42478 11454 42530 11506
rect 6078 11342 6130 11394
rect 6302 11342 6354 11394
rect 6638 11342 6690 11394
rect 8206 11342 8258 11394
rect 8542 11342 8594 11394
rect 8766 11342 8818 11394
rect 14366 11342 14418 11394
rect 14814 11342 14866 11394
rect 15822 11342 15874 11394
rect 16942 11342 16994 11394
rect 21534 11342 21586 11394
rect 26014 11342 26066 11394
rect 31502 11342 31554 11394
rect 31726 11342 31778 11394
rect 41918 11342 41970 11394
rect 42254 11342 42306 11394
rect 4958 11230 5010 11282
rect 5070 11230 5122 11282
rect 5630 11230 5682 11282
rect 8654 11230 8706 11282
rect 9214 11230 9266 11282
rect 9326 11230 9378 11282
rect 11006 11230 11058 11282
rect 14030 11230 14082 11282
rect 15150 11230 15202 11282
rect 15374 11230 15426 11282
rect 26238 11230 26290 11282
rect 31950 11230 32002 11282
rect 32174 11230 32226 11282
rect 32398 11230 32450 11282
rect 32510 11230 32562 11282
rect 38222 11230 38274 11282
rect 42590 11230 42642 11282
rect 48862 11230 48914 11282
rect 52894 11230 52946 11282
rect 53230 11230 53282 11282
rect 5742 11118 5794 11170
rect 6974 11118 7026 11170
rect 8990 11118 9042 11170
rect 11342 11118 11394 11170
rect 14142 11118 14194 11170
rect 15262 11118 15314 11170
rect 16606 11118 16658 11170
rect 24782 11118 24834 11170
rect 36206 11118 36258 11170
rect 40798 11118 40850 11170
rect 48526 11118 48578 11170
rect 49982 11118 50034 11170
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 50558 10950 50610 11002
rect 50662 10950 50714 11002
rect 50766 10950 50818 11002
rect 5070 10782 5122 10834
rect 10894 10782 10946 10834
rect 12014 10782 12066 10834
rect 13246 10782 13298 10834
rect 20750 10782 20802 10834
rect 27358 10782 27410 10834
rect 27918 10782 27970 10834
rect 39454 10782 39506 10834
rect 39902 10782 39954 10834
rect 42702 10782 42754 10834
rect 2494 10670 2546 10722
rect 11678 10670 11730 10722
rect 12798 10670 12850 10722
rect 20974 10670 21026 10722
rect 25230 10670 25282 10722
rect 27246 10670 27298 10722
rect 1822 10558 1874 10610
rect 11006 10558 11058 10610
rect 11454 10558 11506 10610
rect 12126 10558 12178 10610
rect 12574 10558 12626 10610
rect 21086 10558 21138 10610
rect 25566 10558 25618 10610
rect 41022 10558 41074 10610
rect 42814 10558 42866 10610
rect 44270 10558 44322 10610
rect 44494 10558 44546 10610
rect 44830 10558 44882 10610
rect 45726 10558 45778 10610
rect 46398 10558 46450 10610
rect 46622 10558 46674 10610
rect 47182 10558 47234 10610
rect 49198 10558 49250 10610
rect 49422 10558 49474 10610
rect 49646 10558 49698 10610
rect 49758 10558 49810 10610
rect 50318 10558 50370 10610
rect 4622 10446 4674 10498
rect 26014 10446 26066 10498
rect 41582 10446 41634 10498
rect 43262 10446 43314 10498
rect 44382 10446 44434 10498
rect 45278 10446 45330 10498
rect 48974 10446 49026 10498
rect 49310 10446 49362 10498
rect 51102 10446 51154 10498
rect 53230 10446 53282 10498
rect 11118 10334 11170 10386
rect 12238 10334 12290 10386
rect 27358 10334 27410 10386
rect 39230 10334 39282 10386
rect 39902 10334 39954 10386
rect 42702 10334 42754 10386
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 15934 9998 15986 10050
rect 21422 9998 21474 10050
rect 21982 9998 22034 10050
rect 35422 9998 35474 10050
rect 36206 9998 36258 10050
rect 45054 9998 45106 10050
rect 47070 9998 47122 10050
rect 50878 9998 50930 10050
rect 7758 9886 7810 9938
rect 9886 9886 9938 9938
rect 12014 9886 12066 9938
rect 26462 9886 26514 9938
rect 30270 9886 30322 9938
rect 34862 9886 34914 9938
rect 45166 9886 45218 9938
rect 50766 9886 50818 9938
rect 6974 9774 7026 9826
rect 21310 9774 21362 9826
rect 22094 9774 22146 9826
rect 22766 9774 22818 9826
rect 23102 9774 23154 9826
rect 25790 9774 25842 9826
rect 27358 9774 27410 9826
rect 28030 9774 28082 9826
rect 32734 9774 32786 9826
rect 33406 9774 33458 9826
rect 33854 9774 33906 9826
rect 35646 9774 35698 9826
rect 37102 9774 37154 9826
rect 38222 9774 38274 9826
rect 38670 9774 38722 9826
rect 39006 9774 39058 9826
rect 39230 9774 39282 9826
rect 41470 9774 41522 9826
rect 41918 9774 41970 9826
rect 45054 9774 45106 9826
rect 45502 9774 45554 9826
rect 46846 9774 46898 9826
rect 47406 9774 47458 9826
rect 47966 9774 48018 9826
rect 16046 9662 16098 9714
rect 27806 9662 27858 9714
rect 32958 9662 33010 9714
rect 33518 9662 33570 9714
rect 34638 9662 34690 9714
rect 35982 9662 36034 9714
rect 37998 9662 38050 9714
rect 40462 9662 40514 9714
rect 43598 9662 43650 9714
rect 46958 9662 47010 9714
rect 48862 9662 48914 9714
rect 49198 9662 49250 9714
rect 49534 9662 49586 9714
rect 49870 9662 49922 9714
rect 10334 9550 10386 9602
rect 16718 9550 16770 9602
rect 21422 9550 21474 9602
rect 21982 9550 22034 9602
rect 22878 9550 22930 9602
rect 26014 9550 26066 9602
rect 27694 9550 27746 9602
rect 30718 9550 30770 9602
rect 31166 9550 31218 9602
rect 33070 9550 33122 9602
rect 33742 9550 33794 9602
rect 35310 9550 35362 9602
rect 37326 9550 37378 9602
rect 38894 9550 38946 9602
rect 40126 9550 40178 9602
rect 44270 9550 44322 9602
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 50558 9382 50610 9434
rect 50662 9382 50714 9434
rect 50766 9382 50818 9434
rect 7310 9214 7362 9266
rect 7758 9214 7810 9266
rect 13246 9214 13298 9266
rect 25342 9214 25394 9266
rect 31502 9214 31554 9266
rect 35646 9214 35698 9266
rect 35870 9214 35922 9266
rect 37662 9214 37714 9266
rect 42702 9214 42754 9266
rect 46174 9214 46226 9266
rect 46622 9214 46674 9266
rect 52894 9214 52946 9266
rect 4734 9102 4786 9154
rect 10670 9102 10722 9154
rect 14366 9102 14418 9154
rect 25566 9102 25618 9154
rect 27694 9102 27746 9154
rect 35422 9102 35474 9154
rect 4062 8990 4114 9042
rect 9886 8990 9938 9042
rect 13694 8990 13746 9042
rect 17390 8990 17442 9042
rect 25678 8990 25730 9042
rect 27022 8990 27074 9042
rect 30942 8990 30994 9042
rect 39902 8990 39954 9042
rect 40350 8990 40402 9042
rect 41694 8990 41746 9042
rect 43038 8990 43090 9042
rect 45502 8990 45554 9042
rect 45726 8990 45778 9042
rect 49422 8990 49474 9042
rect 53230 8990 53282 9042
rect 6862 8878 6914 8930
rect 7198 8878 7250 8930
rect 12798 8878 12850 8930
rect 13134 8878 13186 8930
rect 16494 8878 16546 8930
rect 18174 8878 18226 8930
rect 20302 8878 20354 8930
rect 26574 8878 26626 8930
rect 29822 8878 29874 8930
rect 30718 8878 30770 8930
rect 35534 8878 35586 8930
rect 41470 8878 41522 8930
rect 45390 8878 45442 8930
rect 48750 8878 48802 8930
rect 49534 8878 49586 8930
rect 52670 8878 52722 8930
rect 30606 8766 30658 8818
rect 39678 8766 39730 8818
rect 41246 8766 41298 8818
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 13582 8318 13634 8370
rect 17054 8318 17106 8370
rect 19406 8318 19458 8370
rect 25902 8318 25954 8370
rect 32398 8318 32450 8370
rect 34526 8318 34578 8370
rect 41470 8318 41522 8370
rect 45390 8318 45442 8370
rect 45838 8318 45890 8370
rect 49310 8318 49362 8370
rect 7870 8206 7922 8258
rect 8542 8206 8594 8258
rect 8990 8206 9042 8258
rect 20078 8206 20130 8258
rect 20526 8206 20578 8258
rect 20750 8206 20802 8258
rect 22206 8206 22258 8258
rect 22654 8206 22706 8258
rect 23102 8206 23154 8258
rect 30494 8206 30546 8258
rect 31278 8206 31330 8258
rect 31614 8206 31666 8258
rect 41022 8206 41074 8258
rect 45166 8206 45218 8258
rect 47742 8206 47794 8258
rect 48862 8206 48914 8258
rect 49086 8206 49138 8258
rect 8654 8094 8706 8146
rect 8878 8094 8930 8146
rect 19742 8094 19794 8146
rect 20414 8094 20466 8146
rect 23774 8094 23826 8146
rect 38334 8094 38386 8146
rect 41806 8094 41858 8146
rect 41918 8094 41970 8146
rect 48078 8094 48130 8146
rect 48638 8094 48690 8146
rect 49534 8094 49586 8146
rect 50542 8094 50594 8146
rect 7982 7982 8034 8034
rect 8094 7982 8146 8034
rect 9550 7982 9602 8034
rect 19518 7982 19570 8034
rect 20302 7982 20354 8034
rect 22094 7982 22146 8034
rect 22318 7982 22370 8034
rect 22430 7982 22482 8034
rect 26350 7982 26402 8034
rect 30158 7982 30210 8034
rect 37998 7982 38050 8034
rect 38222 7982 38274 8034
rect 42142 7982 42194 8034
rect 42478 7982 42530 8034
rect 48190 7982 48242 8034
rect 48414 7982 48466 8034
rect 49646 7982 49698 8034
rect 50654 7982 50706 8034
rect 52670 7982 52722 8034
rect 53006 7982 53058 8034
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 50558 7814 50610 7866
rect 50662 7814 50714 7866
rect 50766 7814 50818 7866
rect 8318 7646 8370 7698
rect 8990 7646 9042 7698
rect 13918 7646 13970 7698
rect 20078 7646 20130 7698
rect 20862 7646 20914 7698
rect 23550 7646 23602 7698
rect 29038 7646 29090 7698
rect 29374 7646 29426 7698
rect 30270 7646 30322 7698
rect 33182 7646 33234 7698
rect 35982 7646 36034 7698
rect 41022 7646 41074 7698
rect 42366 7646 42418 7698
rect 43374 7646 43426 7698
rect 44046 7646 44098 7698
rect 44270 7646 44322 7698
rect 48078 7646 48130 7698
rect 48638 7646 48690 7698
rect 8206 7534 8258 7586
rect 19630 7534 19682 7586
rect 21982 7534 22034 7586
rect 23326 7534 23378 7586
rect 27246 7534 27298 7586
rect 27582 7534 27634 7586
rect 39566 7534 39618 7586
rect 42142 7534 42194 7586
rect 42814 7534 42866 7586
rect 45502 7534 45554 7586
rect 46510 7534 46562 7586
rect 47742 7534 47794 7586
rect 47966 7534 48018 7586
rect 51102 7534 51154 7586
rect 8542 7422 8594 7474
rect 19854 7422 19906 7474
rect 20190 7422 20242 7474
rect 22318 7422 22370 7474
rect 30046 7422 30098 7474
rect 40350 7422 40402 7474
rect 42590 7422 42642 7474
rect 44830 7422 44882 7474
rect 45726 7422 45778 7474
rect 46286 7422 46338 7474
rect 48190 7422 48242 7474
rect 49310 7422 49362 7474
rect 49534 7422 49586 7474
rect 49982 7422 50034 7474
rect 50318 7422 50370 7474
rect 14030 7310 14082 7362
rect 19966 7310 20018 7362
rect 20638 7310 20690 7362
rect 20750 7310 20802 7362
rect 23662 7310 23714 7362
rect 37438 7310 37490 7362
rect 53230 7310 53282 7362
rect 42254 7198 42306 7250
rect 49086 7198 49138 7250
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 26798 6862 26850 6914
rect 37550 6862 37602 6914
rect 37774 6862 37826 6914
rect 38222 6862 38274 6914
rect 42254 6862 42306 6914
rect 42926 6862 42978 6914
rect 49870 6862 49922 6914
rect 53006 6862 53058 6914
rect 8542 6750 8594 6802
rect 18286 6750 18338 6802
rect 32174 6750 32226 6802
rect 35758 6750 35810 6802
rect 36094 6750 36146 6802
rect 36206 6750 36258 6802
rect 38334 6750 38386 6802
rect 38782 6750 38834 6802
rect 42030 6750 42082 6802
rect 46062 6750 46114 6802
rect 50094 6750 50146 6802
rect 53230 6750 53282 6802
rect 7758 6638 7810 6690
rect 11342 6638 11394 6690
rect 15038 6638 15090 6690
rect 15374 6638 15426 6690
rect 16158 6638 16210 6690
rect 25566 6638 25618 6690
rect 27806 6638 27858 6690
rect 29486 6638 29538 6690
rect 32286 6638 32338 6690
rect 32958 6638 33010 6690
rect 36430 6638 36482 6690
rect 38222 6638 38274 6690
rect 42478 6638 42530 6690
rect 46286 6638 46338 6690
rect 49086 6638 49138 6690
rect 49310 6638 49362 6690
rect 49646 6638 49698 6690
rect 50318 6638 50370 6690
rect 51550 6638 51602 6690
rect 51998 6638 52050 6690
rect 25790 6526 25842 6578
rect 26910 6526 26962 6578
rect 27470 6526 27522 6578
rect 31726 6526 31778 6578
rect 31950 6526 32002 6578
rect 33630 6526 33682 6578
rect 39230 6526 39282 6578
rect 41806 6526 41858 6578
rect 45166 6526 45218 6578
rect 45502 6526 45554 6578
rect 46734 6526 46786 6578
rect 47406 6526 47458 6578
rect 52670 6526 52722 6578
rect 10782 6414 10834 6466
rect 26798 6414 26850 6466
rect 27582 6414 27634 6466
rect 29262 6414 29314 6466
rect 32510 6414 32562 6466
rect 49870 6414 49922 6466
rect 51326 6414 51378 6466
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 50558 6246 50610 6298
rect 50662 6246 50714 6298
rect 50766 6246 50818 6298
rect 14702 6078 14754 6130
rect 19742 6078 19794 6130
rect 21646 6078 21698 6130
rect 21758 6078 21810 6130
rect 22430 6078 22482 6130
rect 25566 6078 25618 6130
rect 33070 6078 33122 6130
rect 33294 6078 33346 6130
rect 35870 6078 35922 6130
rect 36878 6078 36930 6130
rect 42702 6078 42754 6130
rect 49198 6078 49250 6130
rect 12126 5966 12178 6018
rect 18958 5966 19010 6018
rect 19966 5966 20018 6018
rect 22878 5966 22930 6018
rect 25230 5966 25282 6018
rect 36206 5966 36258 6018
rect 36318 5966 36370 6018
rect 42030 5966 42082 6018
rect 49870 5966 49922 6018
rect 11342 5854 11394 5906
rect 19630 5854 19682 5906
rect 20190 5854 20242 5906
rect 21310 5854 21362 5906
rect 21422 5854 21474 5906
rect 22206 5854 22258 5906
rect 22654 5854 22706 5906
rect 33742 5854 33794 5906
rect 35982 5854 36034 5906
rect 37214 5854 37266 5906
rect 42366 5854 42418 5906
rect 42590 5854 42642 5906
rect 50318 5854 50370 5906
rect 14254 5742 14306 5794
rect 19854 5742 19906 5794
rect 21534 5742 21586 5794
rect 22542 5742 22594 5794
rect 33182 5742 33234 5794
rect 49534 5742 49586 5794
rect 51102 5742 51154 5794
rect 53230 5742 53282 5794
rect 18846 5630 18898 5682
rect 19182 5630 19234 5682
rect 41806 5630 41858 5682
rect 49982 5630 50034 5682
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19182 5294 19234 5346
rect 22766 5294 22818 5346
rect 31502 5294 31554 5346
rect 38334 5294 38386 5346
rect 45614 5294 45666 5346
rect 15262 5182 15314 5234
rect 17390 5182 17442 5234
rect 18846 5182 18898 5234
rect 22430 5182 22482 5234
rect 29374 5182 29426 5234
rect 29598 5182 29650 5234
rect 30606 5182 30658 5234
rect 36430 5182 36482 5234
rect 40574 5182 40626 5234
rect 44830 5182 44882 5234
rect 46622 5182 46674 5234
rect 47630 5182 47682 5234
rect 48190 5182 48242 5234
rect 14590 5070 14642 5122
rect 17838 5070 17890 5122
rect 25790 5070 25842 5122
rect 26126 5070 26178 5122
rect 27918 5070 27970 5122
rect 28254 5070 28306 5122
rect 28590 5070 28642 5122
rect 29710 5070 29762 5122
rect 30158 5070 30210 5122
rect 31614 5070 31666 5122
rect 37214 5070 37266 5122
rect 37998 5070 38050 5122
rect 38782 5070 38834 5122
rect 46062 5070 46114 5122
rect 46286 5070 46338 5122
rect 48638 5070 48690 5122
rect 49086 5070 49138 5122
rect 18958 4958 19010 5010
rect 22542 4958 22594 5010
rect 28142 4958 28194 5010
rect 28366 4958 28418 5010
rect 29150 4958 29202 5010
rect 38894 4958 38946 5010
rect 46510 4958 46562 5010
rect 24670 4846 24722 4898
rect 26014 4846 26066 4898
rect 29710 4846 29762 4898
rect 37438 4846 37490 4898
rect 39790 4846 39842 4898
rect 44942 4846 44994 4898
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 50558 4678 50610 4730
rect 50662 4678 50714 4730
rect 50766 4678 50818 4730
rect 16830 4510 16882 4562
rect 36094 4510 36146 4562
rect 40238 4510 40290 4562
rect 14926 4398 14978 4450
rect 18174 4398 18226 4450
rect 22318 4398 22370 4450
rect 26014 4398 26066 4450
rect 30046 4398 30098 4450
rect 33854 4398 33906 4450
rect 37662 4398 37714 4450
rect 41694 4398 41746 4450
rect 44942 4398 44994 4450
rect 47854 4398 47906 4450
rect 48190 4398 48242 4450
rect 50878 4398 50930 4450
rect 14366 4286 14418 4338
rect 17390 4286 17442 4338
rect 21646 4286 21698 4338
rect 25230 4286 25282 4338
rect 29262 4286 29314 4338
rect 33070 4286 33122 4338
rect 36990 4286 37042 4338
rect 41022 4286 41074 4338
rect 44270 4286 44322 4338
rect 47518 4286 47570 4338
rect 51662 4286 51714 4338
rect 3614 4174 3666 4226
rect 3726 4174 3778 4226
rect 20302 4174 20354 4226
rect 24446 4174 24498 4226
rect 28142 4174 28194 4226
rect 28814 4174 28866 4226
rect 32174 4174 32226 4226
rect 39790 4174 39842 4226
rect 43822 4174 43874 4226
rect 47070 4174 47122 4226
rect 48750 4174 48802 4226
rect 12126 4062 12178 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 12462 3614 12514 3666
rect 25006 3614 25058 3666
rect 29038 3614 29090 3666
rect 29822 3614 29874 3666
rect 36990 3614 37042 3666
rect 40238 3614 40290 3666
rect 50430 3614 50482 3666
rect 52670 3614 52722 3666
rect 11902 3502 11954 3554
rect 35534 3502 35586 3554
rect 35982 3502 36034 3554
rect 46958 3502 47010 3554
rect 47630 3502 47682 3554
rect 48526 3502 48578 3554
rect 2718 3390 2770 3442
rect 2942 3390 2994 3442
rect 3278 3390 3330 3442
rect 10110 3390 10162 3442
rect 39342 3390 39394 3442
rect 39790 3390 39842 3442
rect 43150 3390 43202 3442
rect 43598 3390 43650 3442
rect 43934 3390 43986 3442
rect 52446 3390 52498 3442
rect 53230 3390 53282 3442
rect 16942 3278 16994 3330
rect 20862 3278 20914 3330
rect 25342 3278 25394 3330
rect 47406 3278 47458 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
rect 50558 3110 50610 3162
rect 50662 3110 50714 3162
rect 50766 3110 50818 3162
<< metal2 >>
rect 13664 54200 13776 55000
rect 41216 54200 41328 55000
rect 4476 50988 4740 50998
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4476 50922 4740 50932
rect 13692 50372 13748 54200
rect 19836 51772 20100 51782
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 19836 51706 20100 51716
rect 41244 51604 41300 54200
rect 50428 51938 50484 51950
rect 50428 51886 50430 51938
rect 50482 51886 50484 51938
rect 41468 51604 41524 51614
rect 41244 51602 41524 51604
rect 41244 51550 41246 51602
rect 41298 51550 41470 51602
rect 41522 51550 41524 51602
rect 41244 51548 41524 51550
rect 50428 51604 50484 51886
rect 51660 51938 51716 51950
rect 51660 51886 51662 51938
rect 51714 51886 51716 51938
rect 50556 51772 50820 51782
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50556 51706 50820 51716
rect 50540 51604 50596 51614
rect 50428 51602 50596 51604
rect 50428 51550 50542 51602
rect 50594 51550 50596 51602
rect 50428 51548 50596 51550
rect 41244 51538 41300 51548
rect 41468 51538 41524 51548
rect 50540 51538 50596 51548
rect 51100 51604 51156 51614
rect 41804 51492 41860 51502
rect 41580 51490 41860 51492
rect 41580 51438 41806 51490
rect 41858 51438 41860 51490
rect 41580 51436 41860 51438
rect 35196 50988 35460 50998
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 41580 50932 41636 51436
rect 41804 51426 41860 51436
rect 35196 50922 35460 50932
rect 40796 50876 41636 50932
rect 49644 51380 49700 51390
rect 18508 50708 18564 50718
rect 31052 50708 31108 50718
rect 18508 50706 18676 50708
rect 18508 50654 18510 50706
rect 18562 50654 18676 50706
rect 18508 50652 18676 50654
rect 18508 50642 18564 50652
rect 13692 50306 13748 50316
rect 15708 50594 15764 50606
rect 15708 50542 15710 50594
rect 15762 50542 15764 50594
rect 13580 49700 13636 49710
rect 4476 49420 4740 49430
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4476 49354 4740 49364
rect 13580 49026 13636 49644
rect 15708 49700 15764 50542
rect 16380 50484 16436 50494
rect 16380 50390 16436 50428
rect 17724 50484 17780 50494
rect 17724 50034 17780 50428
rect 18620 50428 18676 50652
rect 24332 50652 24724 50708
rect 24332 50594 24388 50652
rect 24332 50542 24334 50594
rect 24386 50542 24388 50594
rect 24332 50530 24388 50542
rect 24668 50596 24724 50652
rect 31052 50706 31220 50708
rect 31052 50654 31054 50706
rect 31106 50654 31220 50706
rect 31052 50652 31220 50654
rect 31052 50642 31108 50652
rect 24780 50596 24836 50606
rect 27132 50596 27188 50606
rect 24668 50594 24836 50596
rect 24668 50542 24782 50594
rect 24834 50542 24836 50594
rect 24668 50540 24836 50542
rect 24780 50530 24836 50540
rect 26796 50594 27188 50596
rect 26796 50542 27134 50594
rect 27186 50542 27188 50594
rect 26796 50540 27188 50542
rect 20748 50484 20804 50494
rect 18620 50372 18788 50428
rect 17724 49982 17726 50034
rect 17778 49982 17780 50034
rect 17724 49970 17780 49982
rect 18508 49924 18564 49934
rect 18396 49922 18564 49924
rect 18396 49870 18510 49922
rect 18562 49870 18564 49922
rect 18396 49868 18564 49870
rect 17388 49810 17444 49822
rect 17388 49758 17390 49810
rect 17442 49758 17444 49810
rect 15708 49634 15764 49644
rect 16492 49700 16548 49710
rect 13580 48974 13582 49026
rect 13634 48974 13636 49026
rect 13580 48962 13636 48974
rect 16380 49138 16436 49150
rect 16380 49086 16382 49138
rect 16434 49086 16436 49138
rect 14252 48914 14308 48926
rect 14252 48862 14254 48914
rect 14306 48862 14308 48914
rect 4476 47852 4740 47862
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4476 47786 4740 47796
rect 11340 47460 11396 47470
rect 4476 46284 4740 46294
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4476 46218 4740 46228
rect 8764 45890 8820 45902
rect 8764 45838 8766 45890
rect 8818 45838 8820 45890
rect 4476 44716 4740 44726
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4476 44650 4740 44660
rect 4476 43148 4740 43158
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4476 43082 4740 43092
rect 8764 42756 8820 45838
rect 9436 45778 9492 45790
rect 9436 45726 9438 45778
rect 9490 45726 9492 45778
rect 9436 45332 9492 45726
rect 9436 45266 9492 45276
rect 11340 45106 11396 47404
rect 14028 47460 14084 47470
rect 14028 47366 14084 47404
rect 13244 47348 13300 47358
rect 13244 46898 13300 47292
rect 14140 47348 14196 47358
rect 14140 47254 14196 47292
rect 14252 47234 14308 48862
rect 14588 47460 14644 47470
rect 14588 47458 14756 47460
rect 14588 47406 14590 47458
rect 14642 47406 14756 47458
rect 14588 47404 14756 47406
rect 14588 47394 14644 47404
rect 14252 47182 14254 47234
rect 14306 47182 14308 47234
rect 14252 47170 14308 47182
rect 13244 46846 13246 46898
rect 13298 46846 13300 46898
rect 13244 46834 13300 46846
rect 14700 46898 14756 47404
rect 14700 46846 14702 46898
rect 14754 46846 14756 46898
rect 14700 46834 14756 46846
rect 12012 46788 12068 46798
rect 11676 46786 12068 46788
rect 11676 46734 12014 46786
rect 12066 46734 12068 46786
rect 11676 46732 12068 46734
rect 11564 46002 11620 46014
rect 11564 45950 11566 46002
rect 11618 45950 11620 46002
rect 11564 45556 11620 45950
rect 11564 45490 11620 45500
rect 11564 45332 11620 45342
rect 11564 45238 11620 45276
rect 11340 45054 11342 45106
rect 11394 45054 11396 45106
rect 11228 43764 11284 43774
rect 11340 43764 11396 45054
rect 11564 45108 11620 45118
rect 11676 45108 11732 46732
rect 12012 46722 12068 46732
rect 12236 46788 12292 46798
rect 12236 46694 12292 46732
rect 14028 46788 14084 46798
rect 12348 46676 12404 46686
rect 11900 46562 11956 46574
rect 11900 46510 11902 46562
rect 11954 46510 11956 46562
rect 11788 45220 11844 45230
rect 11788 45126 11844 45164
rect 11564 45106 11732 45108
rect 11564 45054 11566 45106
rect 11618 45054 11732 45106
rect 11564 45052 11732 45054
rect 11564 45042 11620 45052
rect 11564 44098 11620 44110
rect 11564 44046 11566 44098
rect 11618 44046 11620 44098
rect 11564 43764 11620 44046
rect 11228 43762 11396 43764
rect 11228 43710 11230 43762
rect 11282 43710 11396 43762
rect 11228 43708 11396 43710
rect 11228 43698 11284 43708
rect 10892 43540 10948 43550
rect 10780 43484 10892 43540
rect 9660 43428 9716 43438
rect 9660 42866 9716 43372
rect 9660 42814 9662 42866
rect 9714 42814 9716 42866
rect 9660 42802 9716 42814
rect 8876 42756 8932 42766
rect 8764 42754 8932 42756
rect 8764 42702 8878 42754
rect 8930 42702 8932 42754
rect 8764 42700 8932 42702
rect 5068 41970 5124 41982
rect 5068 41918 5070 41970
rect 5122 41918 5124 41970
rect 5068 41860 5124 41918
rect 4476 41580 4740 41590
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4476 41514 4740 41524
rect 4476 40012 4740 40022
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4476 39946 4740 39956
rect 5068 39732 5124 41804
rect 5740 41858 5796 41870
rect 5740 41806 5742 41858
rect 5794 41806 5796 41858
rect 5740 40626 5796 41806
rect 7868 41858 7924 41870
rect 7868 41806 7870 41858
rect 7922 41806 7924 41858
rect 7868 40852 7924 41806
rect 8316 41860 8372 41870
rect 8316 41766 8372 41804
rect 8876 41860 8932 42700
rect 8876 41794 8932 41804
rect 9884 41860 9940 41870
rect 7868 40796 8148 40852
rect 5740 40574 5742 40626
rect 5794 40574 5796 40626
rect 5740 40562 5796 40574
rect 5852 40572 6580 40628
rect 5068 39666 5124 39676
rect 5404 40402 5460 40414
rect 5404 40350 5406 40402
rect 5458 40350 5460 40402
rect 4956 39508 5012 39518
rect 4956 39414 5012 39452
rect 5068 39396 5124 39406
rect 5068 39302 5124 39340
rect 5404 38612 5460 40350
rect 5740 40404 5796 40414
rect 5852 40404 5908 40572
rect 5740 40402 5908 40404
rect 5740 40350 5742 40402
rect 5794 40350 5908 40402
rect 5740 40348 5908 40350
rect 5964 40402 6020 40414
rect 5964 40350 5966 40402
rect 6018 40350 6020 40402
rect 5740 40338 5796 40348
rect 5964 39842 6020 40350
rect 5964 39790 5966 39842
rect 6018 39790 6020 39842
rect 5964 39778 6020 39790
rect 6524 39842 6580 40572
rect 6524 39790 6526 39842
rect 6578 39790 6580 39842
rect 6524 39778 6580 39790
rect 7980 40514 8036 40526
rect 7980 40462 7982 40514
rect 8034 40462 8036 40514
rect 5628 39508 5684 39518
rect 5516 39506 5684 39508
rect 5516 39454 5630 39506
rect 5682 39454 5684 39506
rect 5516 39452 5684 39454
rect 5516 39396 5572 39452
rect 5628 39442 5684 39452
rect 6076 39506 6132 39518
rect 6412 39508 6468 39518
rect 6076 39454 6078 39506
rect 6130 39454 6132 39506
rect 5516 39330 5572 39340
rect 5852 39394 5908 39406
rect 5852 39342 5854 39394
rect 5906 39342 5908 39394
rect 5852 38668 5908 39342
rect 6076 39396 6132 39454
rect 6076 39330 6132 39340
rect 6188 39506 6468 39508
rect 6188 39454 6414 39506
rect 6466 39454 6468 39506
rect 6188 39452 6468 39454
rect 5404 38546 5460 38556
rect 5516 38612 5908 38668
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5516 38052 5572 38612
rect 4620 37996 5012 38052
rect 1820 37266 1876 37278
rect 1820 37214 1822 37266
rect 1874 37214 1876 37266
rect 1820 35924 1876 37214
rect 2492 37156 2548 37166
rect 2492 37062 2548 37100
rect 4620 37154 4676 37996
rect 4956 37938 5012 37996
rect 5180 37996 5572 38052
rect 5628 38332 6020 38388
rect 4956 37886 4958 37938
rect 5010 37886 5012 37938
rect 4956 37874 5012 37886
rect 5068 37938 5124 37950
rect 5068 37886 5070 37938
rect 5122 37886 5124 37938
rect 4732 37828 4788 37838
rect 5068 37828 5124 37886
rect 4732 37826 4900 37828
rect 4732 37774 4734 37826
rect 4786 37774 4900 37826
rect 4732 37772 4900 37774
rect 4732 37762 4788 37772
rect 4844 37266 4900 37772
rect 5068 37762 5124 37772
rect 4844 37214 4846 37266
rect 4898 37214 4900 37266
rect 4844 37202 4900 37214
rect 4620 37102 4622 37154
rect 4674 37102 4676 37154
rect 4620 37044 4676 37102
rect 5068 37156 5124 37166
rect 5068 37062 5124 37100
rect 4620 36978 4676 36988
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 1820 34914 1876 35868
rect 4844 36258 4900 36270
rect 4844 36206 4846 36258
rect 4898 36206 4900 36258
rect 4844 35924 4900 36206
rect 4844 35830 4900 35868
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 5068 35140 5124 35150
rect 1820 34862 1822 34914
rect 1874 34862 1876 34914
rect 1820 32562 1876 34862
rect 4620 35026 4676 35038
rect 4620 34974 4622 35026
rect 4674 34974 4676 35026
rect 4620 34916 4676 34974
rect 5068 34916 5124 35084
rect 4620 34860 5124 34916
rect 2492 34804 2548 34814
rect 2492 34710 2548 34748
rect 5068 34802 5124 34860
rect 5068 34750 5070 34802
rect 5122 34750 5124 34802
rect 4956 34690 5012 34702
rect 4956 34638 4958 34690
rect 5010 34638 5012 34690
rect 4956 34354 5012 34638
rect 5068 34580 5124 34750
rect 5068 34514 5124 34524
rect 5180 34356 5236 37996
rect 5628 37716 5684 38332
rect 5964 38274 6020 38332
rect 5964 38222 5966 38274
rect 6018 38222 6020 38274
rect 5964 38210 6020 38222
rect 5292 37660 5684 37716
rect 5852 38164 5908 38174
rect 5292 37378 5348 37660
rect 5292 37326 5294 37378
rect 5346 37326 5348 37378
rect 5292 37314 5348 37326
rect 5516 37492 5572 37502
rect 5852 37492 5908 38108
rect 6076 38052 6132 38062
rect 5964 37940 6020 37978
rect 6076 37958 6132 37996
rect 5964 37874 6020 37884
rect 6076 37828 6132 37838
rect 6188 37828 6244 39452
rect 6412 39442 6468 39452
rect 6524 39508 6580 39518
rect 7980 39508 8036 40462
rect 8092 40404 8148 40796
rect 8316 40404 8372 40414
rect 8092 40402 8372 40404
rect 8092 40350 8318 40402
rect 8370 40350 8372 40402
rect 8092 40348 8372 40350
rect 8316 39620 8372 40348
rect 8428 39844 8484 39854
rect 8428 39750 8484 39788
rect 9548 39844 9604 39854
rect 9324 39620 9380 39630
rect 8316 39564 8484 39620
rect 8092 39508 8148 39518
rect 7980 39452 8092 39508
rect 6524 39414 6580 39452
rect 7196 39396 7252 39406
rect 6300 39284 6356 39294
rect 6300 38276 6356 39228
rect 7196 39058 7252 39340
rect 7196 39006 7198 39058
rect 7250 39006 7252 39058
rect 7196 38994 7252 39006
rect 7980 39060 8036 39070
rect 7980 38946 8036 39004
rect 7980 38894 7982 38946
rect 8034 38894 8036 38946
rect 7980 38882 8036 38894
rect 8092 38946 8148 39452
rect 8316 39396 8372 39406
rect 8316 39302 8372 39340
rect 8092 38894 8094 38946
rect 8146 38894 8148 38946
rect 8092 38882 8148 38894
rect 8316 39060 8372 39070
rect 7532 38834 7588 38846
rect 7532 38782 7534 38834
rect 7586 38782 7588 38834
rect 7532 38668 7588 38782
rect 8204 38834 8260 38846
rect 8204 38782 8206 38834
rect 8258 38782 8260 38834
rect 8204 38668 8260 38782
rect 6300 38210 6356 38220
rect 6412 38612 6468 38622
rect 6132 37772 6244 37828
rect 5516 37378 5572 37436
rect 5516 37326 5518 37378
rect 5570 37326 5572 37378
rect 5516 37314 5572 37326
rect 5740 37490 5908 37492
rect 5740 37438 5854 37490
rect 5906 37438 5908 37490
rect 5740 37436 5908 37438
rect 5740 36706 5796 37436
rect 5852 37426 5908 37436
rect 5964 37492 6020 37502
rect 6076 37492 6132 37772
rect 6412 37492 6468 38556
rect 7532 38612 8260 38668
rect 5964 37490 6132 37492
rect 5964 37438 5966 37490
rect 6018 37438 6132 37490
rect 5964 37436 6132 37438
rect 6300 37436 6412 37492
rect 5964 37426 6020 37436
rect 6076 37268 6132 37278
rect 6076 37174 6132 37212
rect 5740 36654 5742 36706
rect 5794 36654 5796 36706
rect 5740 36642 5796 36654
rect 5964 36708 6020 36718
rect 5964 36594 6020 36652
rect 5964 36542 5966 36594
rect 6018 36542 6020 36594
rect 5964 36530 6020 36542
rect 6076 36482 6132 36494
rect 6076 36430 6078 36482
rect 6130 36430 6132 36482
rect 6076 36372 6132 36430
rect 6076 36306 6132 36316
rect 5516 35812 5572 35822
rect 5404 35810 5572 35812
rect 5404 35758 5518 35810
rect 5570 35758 5572 35810
rect 5404 35756 5572 35758
rect 5404 35140 5460 35756
rect 5516 35746 5572 35756
rect 5628 35700 5684 35710
rect 5628 35698 6020 35700
rect 5628 35646 5630 35698
rect 5682 35646 6020 35698
rect 5628 35644 6020 35646
rect 5628 35634 5684 35644
rect 5516 35476 5572 35486
rect 5516 35474 5908 35476
rect 5516 35422 5518 35474
rect 5570 35422 5908 35474
rect 5516 35420 5908 35422
rect 5516 35410 5572 35420
rect 5404 35074 5460 35084
rect 5516 34916 5572 34926
rect 4956 34302 4958 34354
rect 5010 34302 5012 34354
rect 4956 34290 5012 34302
rect 5068 34354 5236 34356
rect 5068 34302 5182 34354
rect 5234 34302 5236 34354
rect 5068 34300 5236 34302
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 1820 32510 1822 32562
rect 1874 32510 1876 32562
rect 1820 31948 1876 32510
rect 4620 32900 4676 32910
rect 2492 32452 2548 32462
rect 2492 32358 2548 32396
rect 4620 32450 4676 32844
rect 4620 32398 4622 32450
rect 4674 32398 4676 32450
rect 4620 32386 4676 32398
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 1708 31892 1876 31948
rect 4844 31892 4900 31902
rect 1708 31826 1764 31836
rect 4844 31798 4900 31836
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4956 29988 5012 29998
rect 4844 29932 4956 29988
rect 1820 29426 1876 29438
rect 1820 29374 1822 29426
rect 1874 29374 1876 29426
rect 1820 27074 1876 29374
rect 2492 29314 2548 29326
rect 2492 29262 2494 29314
rect 2546 29262 2548 29314
rect 2492 28866 2548 29262
rect 2492 28814 2494 28866
rect 2546 28814 2548 28866
rect 2492 28802 2548 28814
rect 2828 29316 2884 29326
rect 2828 28866 2884 29260
rect 4620 29314 4676 29326
rect 4620 29262 4622 29314
rect 4674 29262 4676 29314
rect 4620 29204 4676 29262
rect 2828 28814 2830 28866
rect 2882 28814 2884 28866
rect 2828 28802 2884 28814
rect 4284 29148 4620 29204
rect 4284 28868 4340 29148
rect 4620 29138 4676 29148
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 4732 28868 4788 28878
rect 4284 28812 4676 28868
rect 1820 27022 1822 27074
rect 1874 27022 1876 27074
rect 1820 23938 1876 27022
rect 2604 28644 2660 28654
rect 2604 28530 2660 28588
rect 3276 28644 3332 28654
rect 3276 28550 3332 28588
rect 4620 28642 4676 28812
rect 4620 28590 4622 28642
rect 4674 28590 4676 28642
rect 4620 28578 4676 28590
rect 4732 28644 4788 28812
rect 4844 28756 4900 29932
rect 4956 29894 5012 29932
rect 4956 29540 5012 29550
rect 5068 29540 5124 34300
rect 5180 34290 5236 34300
rect 5292 34914 5572 34916
rect 5292 34862 5518 34914
rect 5570 34862 5572 34914
rect 5292 34860 5572 34862
rect 5180 34132 5236 34142
rect 5180 29652 5236 34076
rect 5292 34018 5348 34860
rect 5516 34850 5572 34860
rect 5852 34914 5908 35420
rect 5852 34862 5854 34914
rect 5906 34862 5908 34914
rect 5852 34850 5908 34862
rect 5740 34804 5796 34814
rect 5740 34710 5796 34748
rect 5964 34580 6020 35644
rect 6188 34916 6244 34926
rect 6300 34916 6356 37436
rect 6412 37426 6468 37436
rect 7196 37940 7252 37950
rect 6188 34914 6356 34916
rect 6188 34862 6190 34914
rect 6242 34862 6356 34914
rect 6188 34860 6356 34862
rect 6524 37266 6580 37278
rect 6524 37214 6526 37266
rect 6578 37214 6580 37266
rect 6524 37156 6580 37214
rect 6188 34850 6244 34860
rect 5964 34524 6356 34580
rect 5964 34354 6020 34524
rect 5964 34302 5966 34354
rect 6018 34302 6020 34354
rect 5964 34290 6020 34302
rect 5292 33966 5294 34018
rect 5346 33966 5348 34018
rect 5292 33954 5348 33966
rect 5516 34132 5572 34142
rect 5852 34132 5908 34142
rect 5516 34130 5908 34132
rect 5516 34078 5518 34130
rect 5570 34078 5854 34130
rect 5906 34078 5908 34130
rect 5516 34076 5908 34078
rect 5516 33236 5572 34076
rect 5852 34066 5908 34076
rect 6076 34130 6132 34142
rect 6076 34078 6078 34130
rect 6130 34078 6132 34130
rect 6076 33796 6132 34078
rect 5852 33740 6132 33796
rect 5740 33348 5796 33358
rect 5852 33348 5908 33740
rect 5964 33348 6020 33358
rect 5852 33346 6132 33348
rect 5852 33294 5966 33346
rect 6018 33294 6132 33346
rect 5852 33292 6132 33294
rect 5740 33254 5796 33292
rect 5964 33282 6020 33292
rect 5628 33236 5684 33246
rect 5516 33234 5684 33236
rect 5516 33182 5630 33234
rect 5682 33182 5684 33234
rect 5516 33180 5684 33182
rect 5292 32676 5348 32686
rect 5292 32582 5348 32620
rect 5404 32452 5460 32462
rect 5404 32358 5460 32396
rect 5516 32004 5572 33180
rect 5628 33170 5684 33180
rect 5964 33124 6020 33134
rect 5740 33068 5964 33124
rect 5628 32676 5684 32686
rect 5740 32676 5796 33068
rect 5964 33058 6020 33068
rect 6076 32900 6132 33292
rect 6300 33346 6356 34524
rect 6524 34130 6580 37100
rect 6972 37154 7028 37166
rect 6972 37102 6974 37154
rect 7026 37102 7028 37154
rect 6972 37044 7028 37102
rect 6972 34916 7028 36988
rect 6972 34850 7028 34860
rect 7196 37042 7252 37884
rect 7196 36990 7198 37042
rect 7250 36990 7252 37042
rect 7196 34356 7252 36990
rect 7420 37492 7476 37502
rect 7420 35924 7476 37436
rect 7532 37490 7588 38612
rect 8316 38500 8372 39004
rect 8204 38444 8372 38500
rect 7532 37438 7534 37490
rect 7586 37438 7588 37490
rect 7532 37426 7588 37438
rect 7868 37604 7924 37614
rect 7532 35924 7588 35934
rect 7420 35922 7588 35924
rect 7420 35870 7534 35922
rect 7586 35870 7588 35922
rect 7420 35868 7588 35870
rect 7532 35858 7588 35868
rect 7868 35698 7924 37548
rect 8204 37492 8260 38444
rect 8428 38388 8484 39564
rect 9324 39526 9380 39564
rect 9548 39618 9604 39788
rect 9548 39566 9550 39618
rect 9602 39566 9604 39618
rect 9548 39554 9604 39566
rect 9772 39732 9828 39742
rect 8316 38332 8484 38388
rect 8540 39506 8596 39518
rect 8540 39454 8542 39506
rect 8594 39454 8596 39506
rect 8316 37604 8372 38332
rect 8540 38162 8596 39454
rect 8988 39506 9044 39518
rect 8988 39454 8990 39506
rect 9042 39454 9044 39506
rect 8652 38610 8708 38622
rect 8652 38558 8654 38610
rect 8706 38558 8708 38610
rect 8652 38276 8708 38558
rect 8988 38612 9044 39454
rect 9436 39508 9492 39518
rect 9436 39414 9492 39452
rect 9772 39060 9828 39676
rect 9884 39618 9940 41804
rect 9884 39566 9886 39618
rect 9938 39566 9940 39618
rect 9884 39284 9940 39566
rect 9884 39218 9940 39228
rect 10220 39620 10276 39630
rect 9884 39060 9940 39070
rect 9828 39058 9940 39060
rect 9828 39006 9886 39058
rect 9938 39006 9940 39058
rect 9828 39004 9940 39006
rect 9772 38994 9828 39004
rect 9884 38994 9940 39004
rect 10108 39060 10164 39070
rect 10220 39060 10276 39564
rect 10668 39508 10724 39518
rect 10668 39414 10724 39452
rect 10108 39058 10276 39060
rect 10108 39006 10110 39058
rect 10162 39006 10276 39058
rect 10108 39004 10276 39006
rect 10108 38994 10164 39004
rect 9772 38836 9828 38846
rect 9772 38742 9828 38780
rect 8988 38546 9044 38556
rect 8764 38276 8820 38286
rect 8652 38274 9044 38276
rect 8652 38222 8766 38274
rect 8818 38222 9044 38274
rect 8652 38220 9044 38222
rect 8764 38210 8820 38220
rect 8540 38110 8542 38162
rect 8594 38110 8596 38162
rect 8540 38098 8596 38110
rect 8988 38164 9044 38220
rect 8988 38108 9716 38164
rect 8540 37828 8596 37838
rect 8540 37826 8708 37828
rect 8540 37774 8542 37826
rect 8594 37774 8708 37826
rect 8540 37772 8708 37774
rect 8540 37762 8596 37772
rect 8316 37548 8596 37604
rect 8204 37436 8484 37492
rect 8316 37266 8372 37278
rect 8316 37214 8318 37266
rect 8370 37214 8372 37266
rect 8316 37156 8372 37214
rect 8316 37090 8372 37100
rect 8316 36484 8372 36494
rect 8316 35810 8372 36428
rect 8316 35758 8318 35810
rect 8370 35758 8372 35810
rect 8316 35746 8372 35758
rect 8428 35810 8484 37436
rect 8428 35758 8430 35810
rect 8482 35758 8484 35810
rect 8428 35746 8484 35758
rect 7868 35646 7870 35698
rect 7922 35646 7924 35698
rect 7868 34692 7924 35646
rect 8540 35698 8596 37548
rect 8540 35646 8542 35698
rect 8594 35646 8596 35698
rect 8540 35252 8596 35646
rect 8540 35186 8596 35196
rect 8092 34692 8148 34702
rect 7868 34690 8372 34692
rect 7868 34638 8094 34690
rect 8146 34638 8372 34690
rect 7868 34636 8372 34638
rect 8092 34626 8148 34636
rect 7196 34290 7252 34300
rect 8092 34356 8148 34366
rect 6524 34078 6526 34130
rect 6578 34078 6580 34130
rect 6524 33572 6580 34078
rect 6524 33516 6804 33572
rect 6300 33294 6302 33346
rect 6354 33294 6356 33346
rect 6300 33282 6356 33294
rect 6412 33348 6468 33358
rect 6468 33292 6580 33348
rect 6412 33282 6468 33292
rect 5628 32674 5796 32676
rect 5628 32622 5630 32674
rect 5682 32622 5796 32674
rect 5628 32620 5796 32622
rect 5964 32844 6132 32900
rect 6412 33122 6468 33134
rect 6412 33070 6414 33122
rect 6466 33070 6468 33122
rect 6412 32900 6468 33070
rect 6524 32900 6580 33292
rect 6636 33124 6692 33134
rect 6636 33030 6692 33068
rect 6524 32844 6692 32900
rect 5628 32610 5684 32620
rect 5852 32564 5908 32574
rect 5852 32470 5908 32508
rect 5628 32004 5684 32014
rect 5516 32002 5684 32004
rect 5516 31950 5630 32002
rect 5682 31950 5684 32002
rect 5516 31948 5684 31950
rect 5628 31938 5684 31948
rect 5964 31668 6020 32844
rect 6412 32834 6468 32844
rect 6076 32676 6132 32686
rect 6076 32582 6132 32620
rect 6188 32674 6244 32686
rect 6188 32622 6190 32674
rect 6242 32622 6244 32674
rect 6188 31778 6244 32622
rect 6188 31726 6190 31778
rect 6242 31726 6244 31778
rect 5964 31602 6020 31612
rect 6076 31666 6132 31678
rect 6076 31614 6078 31666
rect 6130 31614 6132 31666
rect 5628 31556 5684 31566
rect 5404 31500 5628 31556
rect 5292 29652 5348 29662
rect 5180 29596 5292 29652
rect 5292 29586 5348 29596
rect 5404 29652 5460 31500
rect 5628 31490 5684 31500
rect 6076 31108 6132 31614
rect 6188 31556 6244 31726
rect 6412 32674 6468 32686
rect 6412 32622 6414 32674
rect 6466 32622 6468 32674
rect 6188 31490 6244 31500
rect 6300 31666 6356 31678
rect 6300 31614 6302 31666
rect 6354 31614 6356 31666
rect 6300 31444 6356 31614
rect 6300 31378 6356 31388
rect 6412 31220 6468 32622
rect 6636 32674 6692 32844
rect 6748 32788 6804 33516
rect 6748 32722 6804 32732
rect 7980 33122 8036 33134
rect 7980 33070 7982 33122
rect 8034 33070 8036 33122
rect 6636 32622 6638 32674
rect 6690 32622 6692 32674
rect 6636 32610 6692 32622
rect 7084 32564 7140 32574
rect 7084 32450 7140 32508
rect 7980 32564 8036 33070
rect 7980 32498 8036 32508
rect 7084 32398 7086 32450
rect 7138 32398 7140 32450
rect 7084 32004 7140 32398
rect 8092 32340 8148 34300
rect 8316 33122 8372 34636
rect 8316 33070 8318 33122
rect 8370 33070 8372 33122
rect 8316 33012 8372 33070
rect 8316 32946 8372 32956
rect 6636 31948 7140 32004
rect 7980 32284 8148 32340
rect 8316 32788 8372 32798
rect 6300 31164 6468 31220
rect 6524 31780 6580 31790
rect 6524 31218 6580 31724
rect 6524 31166 6526 31218
rect 6578 31166 6580 31218
rect 6300 31108 6356 31164
rect 6524 31154 6580 31166
rect 6076 31106 6356 31108
rect 6076 31054 6302 31106
rect 6354 31054 6356 31106
rect 6076 31052 6356 31054
rect 5628 30884 5684 30894
rect 5404 29650 5572 29652
rect 5404 29598 5406 29650
rect 5458 29598 5572 29650
rect 5404 29596 5572 29598
rect 5404 29586 5460 29596
rect 4956 29538 5124 29540
rect 4956 29486 4958 29538
rect 5010 29486 5124 29538
rect 4956 29484 5124 29486
rect 4956 29474 5012 29484
rect 5068 28756 5124 29484
rect 5180 29426 5236 29438
rect 5180 29374 5182 29426
rect 5234 29374 5236 29426
rect 5180 28868 5236 29374
rect 5292 29316 5348 29326
rect 5292 29222 5348 29260
rect 5516 29204 5572 29596
rect 5628 29428 5684 30828
rect 6188 29652 6244 29662
rect 6300 29652 6356 31052
rect 6412 30884 6468 30894
rect 6412 30790 6468 30828
rect 6188 29650 6356 29652
rect 6188 29598 6190 29650
rect 6242 29598 6356 29650
rect 6188 29596 6356 29598
rect 6188 29586 6244 29596
rect 6076 29540 6132 29550
rect 5964 29484 6076 29540
rect 5628 29426 5908 29428
rect 5628 29374 5630 29426
rect 5682 29374 5908 29426
rect 5628 29372 5908 29374
rect 5628 29362 5684 29372
rect 5516 29148 5796 29204
rect 5628 28868 5684 28878
rect 5180 28866 5684 28868
rect 5180 28814 5630 28866
rect 5682 28814 5684 28866
rect 5180 28812 5684 28814
rect 5628 28802 5684 28812
rect 5740 28868 5796 29148
rect 5740 28774 5796 28812
rect 4844 28700 5012 28756
rect 5068 28700 5572 28756
rect 4956 28644 5012 28700
rect 4732 28588 4900 28644
rect 4956 28588 5124 28644
rect 2604 28478 2606 28530
rect 2658 28478 2660 28530
rect 2492 26962 2548 26974
rect 2492 26910 2494 26962
rect 2546 26910 2548 26962
rect 2492 26516 2548 26910
rect 2492 26450 2548 26460
rect 1820 23886 1822 23938
rect 1874 23886 1876 23938
rect 1820 23604 1876 23886
rect 1820 21586 1876 23548
rect 2492 23826 2548 23838
rect 2492 23774 2494 23826
rect 2546 23774 2548 23826
rect 2492 23042 2548 23774
rect 2604 23380 2660 28478
rect 4844 28420 4900 28588
rect 4956 28420 5012 28430
rect 4844 28418 5012 28420
rect 4844 28366 4958 28418
rect 5010 28366 5012 28418
rect 4844 28364 5012 28366
rect 4956 28354 5012 28364
rect 4956 27860 5012 27870
rect 4844 27804 4956 27860
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 4844 27300 4900 27804
rect 4956 27794 5012 27804
rect 4620 27244 4900 27300
rect 4620 27186 4676 27244
rect 4620 27134 4622 27186
rect 4674 27134 4676 27186
rect 4620 27122 4676 27134
rect 5068 27186 5124 28588
rect 5404 27858 5460 27870
rect 5404 27806 5406 27858
rect 5458 27806 5460 27858
rect 5404 27300 5460 27806
rect 5516 27748 5572 28700
rect 5628 27972 5684 27982
rect 5628 27878 5684 27916
rect 5740 27972 5796 27982
rect 5852 27972 5908 29372
rect 5964 28866 6020 29484
rect 6076 29446 6132 29484
rect 6300 29204 6356 29214
rect 5964 28814 5966 28866
rect 6018 28814 6020 28866
rect 5964 28802 6020 28814
rect 6188 29202 6356 29204
rect 6188 29150 6302 29202
rect 6354 29150 6356 29202
rect 6188 29148 6356 29150
rect 6188 28644 6244 29148
rect 6300 29138 6356 29148
rect 5740 27970 5908 27972
rect 5740 27918 5742 27970
rect 5794 27918 5908 27970
rect 5740 27916 5908 27918
rect 6076 28642 6244 28644
rect 6076 28590 6190 28642
rect 6242 28590 6244 28642
rect 6076 28588 6244 28590
rect 5740 27906 5796 27916
rect 5516 27692 5796 27748
rect 5404 27244 5684 27300
rect 5068 27134 5070 27186
rect 5122 27134 5124 27186
rect 5068 26908 5124 27134
rect 5068 26852 5236 26908
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 4396 25396 4452 25406
rect 4284 25340 4396 25396
rect 2828 23716 2884 23726
rect 2604 23378 2772 23380
rect 2604 23326 2606 23378
rect 2658 23326 2772 23378
rect 2604 23324 2772 23326
rect 2604 23314 2660 23324
rect 2492 22990 2494 23042
rect 2546 22990 2548 23042
rect 2492 22978 2548 22990
rect 2716 23044 2772 23324
rect 2828 23266 2884 23660
rect 2828 23214 2830 23266
rect 2882 23214 2884 23266
rect 2828 23202 2884 23214
rect 3276 23044 3332 23054
rect 2716 23042 3332 23044
rect 2716 22990 3278 23042
rect 3330 22990 3332 23042
rect 2716 22988 3332 22990
rect 3276 22978 3332 22988
rect 4284 22596 4340 25340
rect 4396 25330 4452 25340
rect 4732 24836 4788 24846
rect 4788 24780 4900 24836
rect 4732 24742 4788 24780
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4508 24164 4564 24174
rect 4508 23266 4564 24108
rect 4620 24052 4676 24062
rect 4844 24052 4900 24780
rect 5068 24834 5124 24846
rect 5068 24782 5070 24834
rect 5122 24782 5124 24834
rect 5068 24276 5124 24782
rect 4620 24050 4900 24052
rect 4620 23998 4622 24050
rect 4674 23998 4900 24050
rect 4620 23996 4900 23998
rect 4956 24220 5124 24276
rect 5180 24612 5236 26852
rect 5516 26850 5572 26862
rect 5516 26798 5518 26850
rect 5570 26798 5572 26850
rect 5292 26404 5348 26414
rect 5516 26404 5572 26798
rect 5292 26402 5572 26404
rect 5292 26350 5294 26402
rect 5346 26350 5572 26402
rect 5292 26348 5572 26350
rect 5628 26402 5684 27244
rect 5628 26350 5630 26402
rect 5682 26350 5684 26402
rect 5292 26338 5348 26348
rect 5628 26338 5684 26350
rect 5404 26180 5460 26190
rect 5404 26086 5460 26124
rect 5740 25284 5796 27692
rect 5964 27300 6020 27310
rect 6076 27300 6132 28588
rect 6188 28578 6244 28588
rect 5964 27298 6132 27300
rect 5964 27246 5966 27298
rect 6018 27246 6132 27298
rect 5964 27244 6132 27246
rect 6188 28420 6244 28430
rect 6188 27300 6244 28364
rect 5964 26516 6020 27244
rect 6188 27206 6244 27244
rect 6412 27860 6468 27870
rect 6412 27186 6468 27804
rect 6412 27134 6414 27186
rect 6466 27134 6468 27186
rect 6412 27122 6468 27134
rect 5964 26450 6020 26460
rect 5852 26292 5908 26302
rect 6300 26292 6356 26302
rect 6636 26292 6692 31948
rect 7532 31780 7588 31790
rect 6748 31668 6804 31678
rect 6748 31574 6804 31612
rect 7084 31554 7140 31566
rect 7084 31502 7086 31554
rect 7138 31502 7140 31554
rect 6860 31444 6916 31454
rect 6860 30772 6916 31388
rect 7084 31220 7140 31502
rect 7196 31220 7252 31230
rect 7084 31218 7252 31220
rect 7084 31166 7198 31218
rect 7250 31166 7252 31218
rect 7084 31164 7252 31166
rect 6972 30996 7028 31006
rect 6972 30902 7028 30940
rect 7084 30772 7140 30782
rect 6860 30716 7084 30772
rect 7084 29650 7140 30716
rect 7084 29598 7086 29650
rect 7138 29598 7140 29650
rect 7084 29586 7140 29598
rect 6860 29426 6916 29438
rect 6860 29374 6862 29426
rect 6914 29374 6916 29426
rect 6860 29204 6916 29374
rect 6860 29138 6916 29148
rect 6748 27300 6804 27310
rect 6748 26962 6804 27244
rect 6748 26910 6750 26962
rect 6802 26910 6804 26962
rect 6748 26898 6804 26910
rect 7084 27076 7140 27086
rect 7196 27076 7252 31164
rect 7532 31218 7588 31724
rect 7532 31166 7534 31218
rect 7586 31166 7588 31218
rect 7532 31154 7588 31166
rect 7308 29652 7364 29662
rect 7308 29558 7364 29596
rect 7980 29650 8036 32284
rect 7980 29598 7982 29650
rect 8034 29598 8036 29650
rect 7980 29586 8036 29598
rect 8092 30996 8148 31006
rect 7420 29428 7476 29438
rect 7420 29426 7924 29428
rect 7420 29374 7422 29426
rect 7474 29374 7924 29426
rect 7420 29372 7924 29374
rect 7420 29362 7476 29372
rect 7308 29316 7364 29326
rect 7308 28082 7364 29260
rect 7868 29314 7924 29372
rect 7868 29262 7870 29314
rect 7922 29262 7924 29314
rect 7868 29250 7924 29262
rect 7980 29426 8036 29438
rect 7980 29374 7982 29426
rect 8034 29374 8036 29426
rect 7980 28868 8036 29374
rect 7308 28030 7310 28082
rect 7362 28030 7364 28082
rect 7308 28018 7364 28030
rect 7756 28812 8036 28868
rect 7420 27860 7476 27870
rect 7420 27766 7476 27804
rect 7084 27074 7252 27076
rect 7084 27022 7086 27074
rect 7138 27022 7252 27074
rect 7084 27020 7252 27022
rect 7084 26908 7140 27020
rect 5852 26290 6692 26292
rect 5852 26238 5854 26290
rect 5906 26238 6302 26290
rect 6354 26238 6692 26290
rect 5852 26236 6692 26238
rect 5852 26226 5908 26236
rect 6300 26226 6356 26236
rect 6076 25284 6132 25294
rect 5740 25282 6132 25284
rect 5740 25230 6078 25282
rect 6130 25230 6132 25282
rect 5740 25228 6132 25230
rect 5404 24836 5460 24846
rect 5404 24742 5460 24780
rect 4620 23986 4676 23996
rect 4956 23492 5012 24220
rect 5068 24052 5124 24062
rect 5180 24052 5236 24556
rect 6076 24276 6132 25228
rect 6412 25284 6468 25294
rect 6412 25190 6468 25228
rect 6076 24210 6132 24220
rect 6524 24052 6580 24062
rect 5068 24050 5236 24052
rect 5068 23998 5070 24050
rect 5122 23998 5236 24050
rect 5068 23996 5236 23998
rect 5740 24050 6580 24052
rect 5740 23998 6526 24050
rect 6578 23998 6580 24050
rect 5740 23996 6580 23998
rect 5068 23604 5124 23996
rect 5740 23938 5796 23996
rect 6524 23986 6580 23996
rect 5740 23886 5742 23938
rect 5794 23886 5796 23938
rect 5068 23538 5124 23548
rect 5516 23604 5572 23614
rect 4732 23436 4956 23492
rect 4732 23378 4788 23436
rect 4956 23426 5012 23436
rect 5404 23380 5460 23390
rect 4732 23326 4734 23378
rect 4786 23326 4788 23378
rect 4732 23314 4788 23326
rect 5180 23324 5404 23380
rect 4508 23214 4510 23266
rect 4562 23214 4564 23266
rect 4508 23202 4564 23214
rect 4956 23268 5012 23278
rect 4956 23174 5012 23212
rect 5068 22932 5124 22942
rect 5068 22838 5124 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4284 22540 4788 22596
rect 2492 22148 2548 22158
rect 2492 21698 2548 22092
rect 2492 21646 2494 21698
rect 2546 21646 2548 21698
rect 2492 21634 2548 21646
rect 4620 21812 4676 22540
rect 4732 22370 4788 22540
rect 4732 22318 4734 22370
rect 4786 22318 4788 22370
rect 4732 22306 4788 22318
rect 5068 22260 5124 22270
rect 5180 22260 5236 23324
rect 5404 23286 5460 23324
rect 5068 22258 5236 22260
rect 5068 22206 5070 22258
rect 5122 22206 5236 22258
rect 5068 22204 5236 22206
rect 5068 22194 5124 22204
rect 1820 21534 1822 21586
rect 1874 21534 1876 21586
rect 1820 21522 1876 21534
rect 4620 21474 4676 21756
rect 5292 21812 5348 21822
rect 5516 21812 5572 23548
rect 5628 23380 5684 23390
rect 5740 23380 5796 23886
rect 6636 23940 6692 26236
rect 6860 26852 7140 26908
rect 7756 26908 7812 28812
rect 7868 28644 7924 28654
rect 8092 28644 8148 30940
rect 8204 29540 8260 29550
rect 8204 29426 8260 29484
rect 8204 29374 8206 29426
rect 8258 29374 8260 29426
rect 8204 29362 8260 29374
rect 7868 28642 8148 28644
rect 7868 28590 7870 28642
rect 7922 28590 8148 28642
rect 7868 28588 8148 28590
rect 7868 28578 7924 28588
rect 8092 26908 8148 28588
rect 8204 28420 8260 28430
rect 8316 28420 8372 32732
rect 8204 28418 8372 28420
rect 8204 28366 8206 28418
rect 8258 28366 8372 28418
rect 8204 28364 8372 28366
rect 8540 32452 8596 32462
rect 8204 27972 8260 28364
rect 8204 27906 8260 27916
rect 7756 26852 7924 26908
rect 8092 26852 8372 26908
rect 6636 23884 6804 23940
rect 5852 23826 5908 23838
rect 5852 23774 5854 23826
rect 5906 23774 5908 23826
rect 5852 23492 5908 23774
rect 6076 23828 6132 23838
rect 6188 23828 6244 23838
rect 6132 23826 6244 23828
rect 6132 23774 6190 23826
rect 6242 23774 6244 23826
rect 6132 23772 6244 23774
rect 5964 23716 6020 23726
rect 5964 23622 6020 23660
rect 5852 23426 5908 23436
rect 5628 23378 5796 23380
rect 5628 23326 5630 23378
rect 5682 23326 5796 23378
rect 5628 23324 5796 23326
rect 5628 23314 5684 23324
rect 5852 23268 5908 23278
rect 6076 23268 6132 23772
rect 6188 23762 6244 23772
rect 6636 23716 6692 23726
rect 6524 23714 6692 23716
rect 6524 23662 6638 23714
rect 6690 23662 6692 23714
rect 6524 23660 6692 23662
rect 6524 23492 6580 23660
rect 6636 23650 6692 23660
rect 6524 23426 6580 23436
rect 5852 23266 6132 23268
rect 5852 23214 5854 23266
rect 5906 23214 6132 23266
rect 5852 23212 6132 23214
rect 6188 23268 6244 23278
rect 5852 23202 5908 23212
rect 6188 23174 6244 23212
rect 6412 23268 6468 23278
rect 6300 23156 6356 23166
rect 6412 23156 6468 23212
rect 6300 23154 6468 23156
rect 6300 23102 6302 23154
rect 6354 23102 6468 23154
rect 6300 23100 6468 23102
rect 6300 23090 6356 23100
rect 5740 23042 5796 23054
rect 5740 22990 5742 23042
rect 5794 22990 5796 23042
rect 5628 22932 5684 22942
rect 5628 22370 5684 22876
rect 5628 22318 5630 22370
rect 5682 22318 5684 22370
rect 5628 22306 5684 22318
rect 5740 22372 5796 22990
rect 5852 22372 5908 22382
rect 5740 22370 5908 22372
rect 5740 22318 5854 22370
rect 5906 22318 5908 22370
rect 5740 22316 5908 22318
rect 5852 22306 5908 22316
rect 6076 22370 6132 22382
rect 6076 22318 6078 22370
rect 6130 22318 6132 22370
rect 5964 22260 6020 22270
rect 6076 22260 6132 22318
rect 6020 22204 6132 22260
rect 6636 22260 6692 22270
rect 6748 22260 6804 23884
rect 6692 22204 6804 22260
rect 6860 23826 6916 26852
rect 7756 26516 7812 26526
rect 7756 26402 7812 26460
rect 7756 26350 7758 26402
rect 7810 26350 7812 26402
rect 7756 25732 7812 26350
rect 7868 26292 7924 26852
rect 8092 26292 8148 26302
rect 7868 26290 8148 26292
rect 7868 26238 8094 26290
rect 8146 26238 8148 26290
rect 7868 26236 8148 26238
rect 7756 25666 7812 25676
rect 7980 25732 8036 25742
rect 7644 25508 7700 25518
rect 7980 25508 8036 25676
rect 7644 25506 8036 25508
rect 7644 25454 7646 25506
rect 7698 25454 7982 25506
rect 8034 25454 8036 25506
rect 7644 25452 8036 25454
rect 7196 25396 7252 25406
rect 7196 25302 7252 25340
rect 6860 23774 6862 23826
rect 6914 23774 6916 23826
rect 5964 22194 6020 22204
rect 6636 22166 6692 22204
rect 5740 22148 5796 22158
rect 5740 22054 5796 22092
rect 5740 21812 5796 21822
rect 5516 21810 5796 21812
rect 5516 21758 5742 21810
rect 5794 21758 5796 21810
rect 5516 21756 5796 21758
rect 5292 21718 5348 21756
rect 5740 21746 5796 21756
rect 4620 21422 4622 21474
rect 4674 21422 4676 21474
rect 4620 21410 4676 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 6860 20130 6916 23774
rect 7308 25284 7364 25294
rect 7196 23492 7252 23502
rect 7196 23154 7252 23436
rect 7196 23102 7198 23154
rect 7250 23102 7252 23154
rect 7196 23090 7252 23102
rect 7308 21028 7364 25228
rect 7644 24836 7700 25452
rect 7980 25442 8036 25452
rect 8092 25394 8148 26236
rect 8092 25342 8094 25394
rect 8146 25342 8148 25394
rect 8092 25330 8148 25342
rect 8204 25396 8260 25406
rect 8204 25302 8260 25340
rect 7420 24052 7476 24062
rect 7644 24052 7700 24780
rect 7420 24050 7700 24052
rect 7420 23998 7422 24050
rect 7474 23998 7700 24050
rect 7420 23996 7700 23998
rect 7420 23986 7476 23996
rect 7644 23938 7700 23996
rect 7644 23886 7646 23938
rect 7698 23886 7700 23938
rect 7644 23874 7700 23886
rect 8204 23940 8260 23950
rect 8316 23940 8372 26852
rect 8428 26292 8484 26302
rect 8428 25284 8484 26236
rect 8540 25732 8596 32396
rect 8652 31668 8708 37772
rect 8876 37716 8932 37726
rect 8876 37490 8932 37660
rect 8876 37438 8878 37490
rect 8930 37438 8932 37490
rect 8876 37426 8932 37438
rect 8988 37490 9044 38108
rect 9548 37940 9604 37950
rect 8988 37438 8990 37490
rect 9042 37438 9044 37490
rect 8988 37426 9044 37438
rect 9436 37938 9604 37940
rect 9436 37886 9550 37938
rect 9602 37886 9604 37938
rect 9436 37884 9604 37886
rect 8764 37268 8820 37278
rect 8764 37174 8820 37212
rect 9324 37268 9380 37278
rect 9100 36372 9156 36382
rect 9156 36316 9268 36372
rect 9100 36278 9156 36316
rect 8988 35476 9044 35486
rect 8876 35474 9044 35476
rect 8876 35422 8990 35474
rect 9042 35422 9044 35474
rect 8876 35420 9044 35422
rect 8764 34916 8820 34926
rect 8876 34916 8932 35420
rect 8988 35410 9044 35420
rect 8764 34914 8932 34916
rect 8764 34862 8766 34914
rect 8818 34862 8932 34914
rect 8764 34860 8932 34862
rect 8764 34850 8820 34860
rect 8988 34802 9044 34814
rect 8988 34750 8990 34802
rect 9042 34750 9044 34802
rect 8876 34356 8932 34366
rect 8988 34356 9044 34750
rect 8932 34300 9044 34356
rect 8876 34290 8932 34300
rect 9212 33572 9268 36316
rect 8988 33570 9268 33572
rect 8988 33518 9214 33570
rect 9266 33518 9268 33570
rect 8988 33516 9268 33518
rect 8764 33122 8820 33134
rect 8764 33070 8766 33122
rect 8818 33070 8820 33122
rect 8764 33012 8820 33070
rect 8764 32946 8820 32956
rect 8876 32900 8932 32910
rect 8876 31780 8932 32844
rect 8652 30436 8708 31612
rect 8652 30370 8708 30380
rect 8764 31724 8932 31780
rect 8764 26908 8820 31724
rect 8876 31554 8932 31566
rect 8876 31502 8878 31554
rect 8930 31502 8932 31554
rect 8876 30996 8932 31502
rect 8876 30930 8932 30940
rect 8988 28420 9044 33516
rect 9212 33506 9268 33516
rect 9324 32228 9380 37212
rect 9436 36706 9492 37884
rect 9548 37874 9604 37884
rect 9660 37938 9716 38108
rect 9660 37886 9662 37938
rect 9714 37886 9716 37938
rect 9660 37874 9716 37886
rect 9884 37828 9940 37838
rect 9884 37734 9940 37772
rect 10444 37828 10500 37838
rect 9548 37716 9604 37726
rect 9548 37378 9604 37660
rect 9548 37326 9550 37378
rect 9602 37326 9604 37378
rect 9548 37314 9604 37326
rect 9660 37378 9716 37390
rect 9660 37326 9662 37378
rect 9714 37326 9716 37378
rect 9660 37044 9716 37326
rect 9884 37378 9940 37390
rect 9884 37326 9886 37378
rect 9938 37326 9940 37378
rect 9884 37268 9940 37326
rect 10444 37378 10500 37772
rect 10780 37604 10836 43484
rect 10892 43446 10948 43484
rect 11340 43316 11396 43708
rect 11452 43708 11620 43764
rect 11452 43540 11508 43708
rect 11788 43652 11844 43662
rect 11788 43558 11844 43596
rect 11452 43474 11508 43484
rect 11564 43538 11620 43550
rect 11564 43486 11566 43538
rect 11618 43486 11620 43538
rect 11564 43316 11620 43486
rect 11340 43260 11620 43316
rect 11900 42980 11956 46510
rect 12012 45892 12068 45902
rect 12348 45892 12404 46620
rect 13132 46676 13188 46686
rect 12796 46564 12852 46574
rect 12796 46470 12852 46508
rect 13132 46004 13188 46620
rect 13132 45938 13188 45948
rect 13356 46674 13412 46686
rect 13356 46622 13358 46674
rect 13410 46622 13412 46674
rect 13356 46564 13412 46622
rect 13804 46676 13860 46686
rect 13804 46674 13972 46676
rect 13804 46622 13806 46674
rect 13858 46622 13972 46674
rect 13804 46620 13972 46622
rect 13804 46610 13860 46620
rect 12012 45890 12404 45892
rect 12012 45838 12014 45890
rect 12066 45838 12404 45890
rect 12012 45836 12404 45838
rect 12012 45826 12068 45836
rect 12124 45666 12180 45678
rect 12124 45614 12126 45666
rect 12178 45614 12180 45666
rect 12124 45220 12180 45614
rect 12236 45666 12292 45678
rect 12236 45614 12238 45666
rect 12290 45614 12292 45666
rect 12236 45444 12292 45614
rect 12460 45668 12516 45678
rect 13356 45668 13412 46508
rect 13580 45668 13636 45678
rect 13356 45666 13636 45668
rect 13356 45614 13582 45666
rect 13634 45614 13636 45666
rect 13356 45612 13636 45614
rect 12236 45378 12292 45388
rect 12348 45556 12404 45566
rect 12124 45154 12180 45164
rect 12236 45108 12292 45118
rect 12348 45108 12404 45500
rect 12460 45330 12516 45612
rect 13580 45444 13636 45612
rect 13580 45378 13636 45388
rect 13916 45556 13972 46620
rect 14028 45892 14084 46732
rect 14252 46676 14308 46686
rect 14028 45798 14084 45836
rect 14140 46674 14308 46676
rect 14140 46622 14254 46674
rect 14306 46622 14308 46674
rect 14140 46620 14308 46622
rect 12460 45278 12462 45330
rect 12514 45278 12516 45330
rect 12460 45266 12516 45278
rect 12236 45106 12404 45108
rect 12236 45054 12238 45106
rect 12290 45054 12404 45106
rect 12236 45052 12404 45054
rect 13916 45108 13972 45500
rect 14028 45108 14084 45118
rect 13916 45106 14084 45108
rect 13916 45054 14030 45106
rect 14082 45054 14084 45106
rect 13916 45052 14084 45054
rect 12236 43876 12292 45052
rect 14028 45042 14084 45052
rect 14140 45108 14196 46620
rect 14252 46610 14308 46620
rect 14476 46674 14532 46686
rect 14476 46622 14478 46674
rect 14530 46622 14532 46674
rect 14252 46004 14308 46014
rect 14252 45910 14308 45948
rect 14476 45780 14532 46622
rect 14700 46676 14756 46686
rect 15036 46676 15092 46686
rect 14700 46674 15092 46676
rect 14700 46622 14702 46674
rect 14754 46622 15038 46674
rect 15090 46622 15092 46674
rect 14700 46620 15092 46622
rect 14700 46610 14756 46620
rect 15036 46610 15092 46620
rect 15148 46562 15204 46574
rect 15148 46510 15150 46562
rect 15202 46510 15204 46562
rect 14252 45778 14532 45780
rect 14252 45726 14478 45778
rect 14530 45726 14532 45778
rect 14252 45724 14532 45726
rect 14252 45668 14308 45724
rect 14476 45714 14532 45724
rect 14588 45892 14644 45902
rect 14252 45218 14308 45612
rect 14252 45166 14254 45218
rect 14306 45166 14308 45218
rect 14252 45154 14308 45166
rect 14364 45220 14420 45230
rect 14588 45220 14644 45836
rect 14364 45218 14644 45220
rect 14364 45166 14366 45218
rect 14418 45166 14644 45218
rect 14364 45164 14644 45166
rect 15036 45890 15092 45902
rect 15036 45838 15038 45890
rect 15090 45838 15092 45890
rect 14364 45154 14420 45164
rect 12236 43820 12964 43876
rect 12348 43650 12404 43662
rect 12348 43598 12350 43650
rect 12402 43598 12404 43650
rect 12236 43540 12292 43550
rect 12348 43540 12404 43598
rect 12236 43538 12404 43540
rect 12236 43486 12238 43538
rect 12290 43486 12404 43538
rect 12236 43484 12404 43486
rect 12572 43650 12628 43662
rect 12572 43598 12574 43650
rect 12626 43598 12628 43650
rect 12236 43474 12292 43484
rect 12012 43428 12068 43438
rect 12012 43334 12068 43372
rect 11900 42924 12292 42980
rect 11788 42866 11844 42878
rect 11788 42814 11790 42866
rect 11842 42814 11844 42866
rect 11788 42084 11844 42814
rect 12236 42868 12292 42924
rect 12236 42774 12292 42812
rect 12572 42644 12628 43598
rect 12684 43538 12740 43550
rect 12684 43486 12686 43538
rect 12738 43486 12740 43538
rect 12684 43316 12740 43486
rect 12684 43250 12740 43260
rect 12572 42196 12628 42588
rect 12684 42196 12740 42206
rect 12572 42194 12740 42196
rect 12572 42142 12686 42194
rect 12738 42142 12740 42194
rect 12572 42140 12740 42142
rect 12684 42130 12740 42140
rect 11788 42028 12404 42084
rect 12348 41970 12404 42028
rect 12348 41918 12350 41970
rect 12402 41918 12404 41970
rect 12348 40292 12404 41918
rect 12460 40292 12516 40302
rect 12348 40236 12460 40292
rect 12460 40226 12516 40236
rect 12796 39732 12852 39742
rect 12796 39638 12852 39676
rect 10780 37538 10836 37548
rect 11004 39284 11060 39294
rect 10444 37326 10446 37378
rect 10498 37326 10500 37378
rect 10444 37314 10500 37326
rect 9996 37268 10052 37278
rect 9884 37266 10052 37268
rect 9884 37214 9998 37266
rect 10050 37214 10052 37266
rect 9884 37212 10052 37214
rect 9996 37202 10052 37212
rect 10220 37268 10276 37278
rect 10220 37174 10276 37212
rect 10668 37266 10724 37278
rect 10668 37214 10670 37266
rect 10722 37214 10724 37266
rect 9436 36654 9438 36706
rect 9490 36654 9492 36706
rect 9436 36642 9492 36654
rect 9548 36988 9660 37044
rect 9436 36484 9492 36494
rect 9548 36484 9604 36988
rect 9660 36978 9716 36988
rect 9492 36428 9604 36484
rect 9436 36390 9492 36428
rect 10668 36260 10724 37214
rect 11004 37266 11060 39228
rect 11004 37214 11006 37266
rect 11058 37214 11060 37266
rect 11004 37156 11060 37214
rect 11788 37268 11844 37278
rect 11788 37174 11844 37212
rect 10892 36260 10948 36270
rect 10668 36258 10948 36260
rect 10668 36206 10894 36258
rect 10946 36206 10948 36258
rect 10668 36204 10948 36206
rect 10892 35924 10948 36204
rect 10892 35858 10948 35868
rect 11004 35308 11060 37100
rect 12908 36484 12964 43820
rect 14028 43652 14084 43662
rect 14028 43558 14084 43596
rect 14140 43650 14196 45052
rect 15036 44996 15092 45838
rect 15148 45556 15204 46510
rect 15932 45890 15988 45902
rect 15932 45838 15934 45890
rect 15986 45838 15988 45890
rect 15932 45668 15988 45838
rect 15932 45602 15988 45612
rect 15148 45490 15204 45500
rect 16380 45556 16436 49086
rect 16380 45490 16436 45500
rect 16492 48804 16548 49644
rect 16828 48804 16884 48814
rect 16492 48802 16884 48804
rect 16492 48750 16830 48802
rect 16882 48750 16884 48802
rect 16492 48748 16884 48750
rect 16492 45668 16548 48748
rect 16828 48738 16884 48748
rect 17388 47460 17444 49758
rect 17724 49812 17780 49822
rect 18060 49812 18116 49822
rect 17724 49810 17892 49812
rect 17724 49758 17726 49810
rect 17778 49758 17892 49810
rect 17724 49756 17892 49758
rect 17724 49746 17780 49756
rect 17836 49364 17892 49756
rect 18060 49718 18116 49756
rect 17836 49308 18228 49364
rect 18172 49026 18228 49308
rect 18172 48974 18174 49026
rect 18226 48974 18228 49026
rect 18172 48962 18228 48974
rect 18396 48916 18452 49868
rect 18508 49858 18564 49868
rect 18732 49810 18788 50372
rect 18732 49758 18734 49810
rect 18786 49758 18788 49810
rect 18396 48822 18452 48860
rect 18508 48914 18564 48926
rect 18508 48862 18510 48914
rect 18562 48862 18564 48914
rect 18508 48468 18564 48862
rect 18508 48402 18564 48412
rect 17388 47394 17444 47404
rect 18732 46228 18788 49758
rect 18956 50370 19012 50382
rect 18956 50318 18958 50370
rect 19010 50318 19012 50370
rect 18956 49700 19012 50318
rect 19836 50204 20100 50214
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 19836 50138 20100 50148
rect 20748 49922 20804 50428
rect 23996 50482 24052 50494
rect 23996 50430 23998 50482
rect 24050 50430 24052 50482
rect 20748 49870 20750 49922
rect 20802 49870 20804 49922
rect 20748 49858 20804 49870
rect 22764 50372 22820 50382
rect 18956 49634 19012 49644
rect 19292 49812 19348 49822
rect 19292 49250 19348 49756
rect 20076 49810 20132 49822
rect 20076 49758 20078 49810
rect 20130 49758 20132 49810
rect 19628 49700 19684 49710
rect 19628 49606 19684 49644
rect 20076 49700 20132 49758
rect 20076 49634 20132 49644
rect 19292 49198 19294 49250
rect 19346 49198 19348 49250
rect 19292 49186 19348 49198
rect 19964 49084 20468 49140
rect 19628 49028 19684 49038
rect 19628 48934 19684 48972
rect 19964 49026 20020 49084
rect 19964 48974 19966 49026
rect 20018 48974 20020 49026
rect 19964 48962 20020 48974
rect 19516 48916 19572 48926
rect 19404 48804 19460 48814
rect 19404 48710 19460 48748
rect 19516 48356 19572 48860
rect 20300 48916 20356 48926
rect 20300 48822 20356 48860
rect 20188 48804 20244 48814
rect 20188 48710 20244 48748
rect 19836 48636 20100 48646
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 19836 48570 20100 48580
rect 20076 48356 20132 48366
rect 20412 48356 20468 49084
rect 19516 48300 19684 48356
rect 19404 48244 19460 48254
rect 19404 48132 19460 48188
rect 19516 48132 19572 48142
rect 19404 48130 19572 48132
rect 19404 48078 19518 48130
rect 19570 48078 19572 48130
rect 19404 48076 19572 48078
rect 19292 48020 19348 48030
rect 19292 47458 19348 47964
rect 19292 47406 19294 47458
rect 19346 47406 19348 47458
rect 19292 47394 19348 47406
rect 19404 47346 19460 48076
rect 19516 48066 19572 48076
rect 19404 47294 19406 47346
rect 19458 47294 19460 47346
rect 18732 46162 18788 46172
rect 18844 47234 18900 47246
rect 18844 47182 18846 47234
rect 18898 47182 18900 47234
rect 18732 46002 18788 46014
rect 18732 45950 18734 46002
rect 18786 45950 18788 46002
rect 16268 45444 16324 45454
rect 15372 44996 15428 45006
rect 15036 44940 15372 44996
rect 15372 44902 15428 44940
rect 14812 44882 14868 44894
rect 14812 44830 14814 44882
rect 14866 44830 14868 44882
rect 14140 43598 14142 43650
rect 14194 43598 14196 43650
rect 14140 43586 14196 43598
rect 14476 44212 14532 44222
rect 14364 43538 14420 43550
rect 14364 43486 14366 43538
rect 14418 43486 14420 43538
rect 14028 43092 14084 43102
rect 14028 42978 14084 43036
rect 14028 42926 14030 42978
rect 14082 42926 14084 42978
rect 14028 42914 14084 42926
rect 14364 42978 14420 43486
rect 14364 42926 14366 42978
rect 14418 42926 14420 42978
rect 14364 42914 14420 42926
rect 13020 42868 13076 42878
rect 13020 39058 13076 42812
rect 13804 42644 13860 42654
rect 14476 42644 14532 44156
rect 14700 43538 14756 43550
rect 14700 43486 14702 43538
rect 14754 43486 14756 43538
rect 13860 42588 13972 42644
rect 13804 42550 13860 42588
rect 13916 42196 13972 42588
rect 14140 42196 14196 42206
rect 13916 42140 14140 42196
rect 14140 42102 14196 42140
rect 14364 42196 14420 42206
rect 14476 42196 14532 42588
rect 14364 42194 14532 42196
rect 14364 42142 14366 42194
rect 14418 42142 14532 42194
rect 14364 42140 14532 42142
rect 14588 43092 14644 43102
rect 14364 42130 14420 42140
rect 14588 42084 14644 43036
rect 14700 42868 14756 43486
rect 14812 43092 14868 44830
rect 14812 43026 14868 43036
rect 16156 44324 16212 44334
rect 15260 42980 15316 42990
rect 15260 42978 16100 42980
rect 15260 42926 15262 42978
rect 15314 42926 16100 42978
rect 15260 42924 16100 42926
rect 15260 42914 15316 42924
rect 16044 42868 16100 42924
rect 16156 42868 16212 44268
rect 16268 44212 16324 45388
rect 16380 44212 16436 44222
rect 16268 44210 16436 44212
rect 16268 44158 16382 44210
rect 16434 44158 16436 44210
rect 16268 44156 16436 44158
rect 14700 42812 15092 42868
rect 14700 42754 14756 42812
rect 14700 42702 14702 42754
rect 14754 42702 14756 42754
rect 14700 42690 14756 42702
rect 14924 42644 14980 42654
rect 14924 42550 14980 42588
rect 15036 42420 15092 42812
rect 16044 42866 16212 42868
rect 16044 42814 16046 42866
rect 16098 42814 16212 42866
rect 16044 42812 16212 42814
rect 16044 42802 16100 42812
rect 15372 42754 15428 42766
rect 15372 42702 15374 42754
rect 15426 42702 15428 42754
rect 15148 42532 15204 42542
rect 15148 42438 15204 42476
rect 14924 42364 15092 42420
rect 14588 41990 14644 42028
rect 14812 42308 14868 42318
rect 14476 41748 14532 41758
rect 14364 41746 14532 41748
rect 14364 41694 14478 41746
rect 14530 41694 14532 41746
rect 14364 41692 14532 41694
rect 14364 41186 14420 41692
rect 14476 41682 14532 41692
rect 14812 41410 14868 42252
rect 14924 41748 14980 42364
rect 15036 42196 15092 42206
rect 15036 42102 15092 42140
rect 15148 42084 15204 42094
rect 15148 41990 15204 42028
rect 15036 41748 15092 41758
rect 14924 41746 15092 41748
rect 14924 41694 15038 41746
rect 15090 41694 15092 41746
rect 14924 41692 15092 41694
rect 15036 41682 15092 41692
rect 14812 41358 14814 41410
rect 14866 41358 14868 41410
rect 14812 41346 14868 41358
rect 14364 41134 14366 41186
rect 14418 41134 14420 41186
rect 14364 41122 14420 41134
rect 14700 41188 14756 41198
rect 14700 41094 14756 41132
rect 15148 41186 15204 41198
rect 15148 41134 15150 41186
rect 15202 41134 15204 41186
rect 14476 40964 14532 40974
rect 14252 40962 14532 40964
rect 14252 40910 14478 40962
rect 14530 40910 14532 40962
rect 14252 40908 14532 40910
rect 14252 39730 14308 40908
rect 14476 40898 14532 40908
rect 15148 40964 15204 41134
rect 15148 40898 15204 40908
rect 15372 41188 15428 42702
rect 16380 41972 16436 44156
rect 16380 41906 16436 41916
rect 15372 40626 15428 41132
rect 16380 41188 16436 41198
rect 16492 41188 16548 45612
rect 16604 45778 16660 45790
rect 16604 45726 16606 45778
rect 16658 45726 16660 45778
rect 16604 44548 16660 45726
rect 16604 44482 16660 44492
rect 16940 45556 16996 45566
rect 16828 44324 16884 44334
rect 16828 44230 16884 44268
rect 16380 41186 16548 41188
rect 16380 41134 16382 41186
rect 16434 41134 16548 41186
rect 16380 41132 16548 41134
rect 15596 40964 15652 40974
rect 15652 40908 15764 40964
rect 15596 40870 15652 40908
rect 15372 40574 15374 40626
rect 15426 40574 15428 40626
rect 15372 40562 15428 40574
rect 15260 40292 15316 40302
rect 14252 39678 14254 39730
rect 14306 39678 14308 39730
rect 14252 39666 14308 39678
rect 15148 39732 15204 39742
rect 13580 39620 13636 39630
rect 13580 39526 13636 39564
rect 13020 39006 13022 39058
rect 13074 39006 13076 39058
rect 13020 38668 13076 39006
rect 13020 38612 13524 38668
rect 13468 37156 13524 38612
rect 13468 37090 13524 37100
rect 13916 37154 13972 37166
rect 13916 37102 13918 37154
rect 13970 37102 13972 37154
rect 13916 37044 13972 37102
rect 14364 37156 14420 37166
rect 14364 37062 14420 37100
rect 13916 36978 13972 36988
rect 12908 36418 12964 36428
rect 15148 36482 15204 39676
rect 15260 37266 15316 40236
rect 15484 40290 15540 40302
rect 15484 40238 15486 40290
rect 15538 40238 15540 40290
rect 15484 39732 15540 40238
rect 15484 39666 15540 39676
rect 15708 38668 15764 40908
rect 16380 40404 16436 41132
rect 16604 40404 16660 40414
rect 16716 40404 16772 40414
rect 16380 40402 16716 40404
rect 16380 40350 16606 40402
rect 16658 40350 16716 40402
rect 16380 40348 16716 40350
rect 16604 40338 16660 40348
rect 16380 39732 16436 39742
rect 16380 38834 16436 39676
rect 16716 39620 16772 40348
rect 16940 39620 16996 45500
rect 18620 45332 18676 45342
rect 18732 45332 18788 45950
rect 18844 45556 18900 47182
rect 18956 46674 19012 46686
rect 18956 46622 18958 46674
rect 19010 46622 19012 46674
rect 18956 46114 19012 46622
rect 19404 46676 19460 47294
rect 19628 47458 19684 48300
rect 20076 48354 20412 48356
rect 20076 48302 20078 48354
rect 20130 48302 20412 48354
rect 20076 48300 20412 48302
rect 20076 48290 20132 48300
rect 20412 48262 20468 48300
rect 20636 48580 20692 48590
rect 20636 48354 20692 48524
rect 21532 48468 21588 48478
rect 21532 48374 21588 48412
rect 22204 48468 22260 48478
rect 22204 48374 22260 48412
rect 20636 48302 20638 48354
rect 20690 48302 20692 48354
rect 19740 48020 19796 48030
rect 19740 47926 19796 47964
rect 19628 47406 19630 47458
rect 19682 47406 19684 47458
rect 19628 46900 19684 47406
rect 20636 47124 20692 48302
rect 22092 48356 22148 48366
rect 22092 48262 22148 48300
rect 22316 48356 22372 48366
rect 22316 48262 22372 48300
rect 21084 48242 21140 48254
rect 21084 48190 21086 48242
rect 21138 48190 21140 48242
rect 20748 48132 20804 48142
rect 21084 48132 21140 48190
rect 20748 48130 21140 48132
rect 20748 48078 20750 48130
rect 20802 48078 21140 48130
rect 20748 48076 21140 48078
rect 21308 48242 21364 48254
rect 21308 48190 21310 48242
rect 21362 48190 21364 48242
rect 20748 48066 20804 48076
rect 21308 48020 21364 48190
rect 21644 48244 21700 48254
rect 21644 48150 21700 48188
rect 22652 48244 22708 48254
rect 22652 48150 22708 48188
rect 21420 48132 21476 48142
rect 21420 48038 21476 48076
rect 21308 47348 21364 47964
rect 21308 47292 21924 47348
rect 19836 47068 20100 47078
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 19836 47002 20100 47012
rect 20188 47068 20692 47124
rect 19628 46844 20132 46900
rect 20076 46786 20132 46844
rect 20076 46734 20078 46786
rect 20130 46734 20132 46786
rect 20076 46722 20132 46734
rect 19404 46610 19460 46620
rect 19628 46674 19684 46686
rect 19628 46622 19630 46674
rect 19682 46622 19684 46674
rect 18956 46062 18958 46114
rect 19010 46062 19012 46114
rect 18956 46050 19012 46062
rect 19292 46114 19348 46126
rect 19292 46062 19294 46114
rect 19346 46062 19348 46114
rect 19180 45668 19236 45678
rect 19180 45574 19236 45612
rect 18844 45500 19012 45556
rect 18676 45276 18788 45332
rect 18060 45220 18116 45230
rect 18060 45126 18116 45164
rect 18620 45218 18676 45276
rect 18620 45166 18622 45218
rect 18674 45166 18676 45218
rect 18620 45154 18676 45166
rect 18844 45220 18900 45230
rect 18284 45108 18340 45118
rect 18844 45108 18900 45164
rect 18956 45108 19012 45500
rect 19068 45220 19124 45230
rect 19068 45126 19124 45164
rect 18844 45106 19012 45108
rect 18844 45054 18958 45106
rect 19010 45054 19012 45106
rect 18844 45052 19012 45054
rect 18284 45014 18340 45052
rect 18956 45042 19012 45052
rect 18172 44994 18228 45006
rect 18172 44942 18174 44994
rect 18226 44942 18228 44994
rect 18172 44660 18228 44942
rect 19068 44884 19124 44894
rect 18844 44828 19068 44884
rect 17612 44604 18228 44660
rect 18284 44660 18340 44670
rect 17276 44548 17332 44558
rect 17276 44454 17332 44492
rect 17612 44546 17668 44604
rect 18284 44548 18340 44604
rect 17612 44494 17614 44546
rect 17666 44494 17668 44546
rect 17612 44482 17668 44494
rect 18172 44492 18340 44548
rect 17724 44436 17780 44446
rect 17724 44342 17780 44380
rect 17388 44324 17444 44334
rect 18172 44324 18228 44492
rect 18396 44436 18452 44446
rect 17388 44322 17668 44324
rect 17388 44270 17390 44322
rect 17442 44270 17668 44322
rect 17388 44268 17668 44270
rect 17388 44258 17444 44268
rect 17612 43876 17668 44268
rect 18172 44230 18228 44268
rect 18284 44380 18396 44436
rect 17612 43820 18116 43876
rect 18060 43762 18116 43820
rect 18060 43710 18062 43762
rect 18114 43710 18116 43762
rect 17052 43428 17108 43438
rect 17052 41298 17108 43372
rect 18060 41412 18116 43710
rect 18284 43538 18340 44380
rect 18396 44370 18452 44380
rect 18620 44436 18676 44446
rect 18620 44342 18676 44380
rect 18844 44322 18900 44828
rect 19068 44790 19124 44828
rect 18844 44270 18846 44322
rect 18898 44270 18900 44322
rect 18844 44258 18900 44270
rect 19292 44436 19348 46062
rect 19628 45332 19684 46622
rect 20188 46564 20244 47068
rect 21084 46900 21140 46910
rect 21084 46806 21140 46844
rect 20412 46788 20468 46798
rect 20412 46694 20468 46732
rect 20972 46788 21028 46798
rect 20972 46694 21028 46732
rect 20300 46676 20356 46686
rect 20300 46582 20356 46620
rect 20076 46508 20244 46564
rect 20076 45668 20132 46508
rect 21868 46114 21924 47292
rect 21868 46062 21870 46114
rect 21922 46062 21924 46114
rect 21868 46050 21924 46062
rect 22540 46674 22596 46686
rect 22540 46622 22542 46674
rect 22594 46622 22596 46674
rect 22540 46564 22596 46622
rect 22540 46002 22596 46508
rect 22540 45950 22542 46002
rect 22594 45950 22596 46002
rect 22540 45938 22596 45950
rect 22428 45892 22484 45902
rect 22428 45798 22484 45836
rect 22652 45890 22708 45902
rect 22652 45838 22654 45890
rect 22706 45838 22708 45890
rect 20076 45612 20244 45668
rect 19836 45500 20100 45510
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 19836 45434 20100 45444
rect 20188 45332 20244 45612
rect 22652 45556 22708 45838
rect 19628 45266 19684 45276
rect 20076 45276 20244 45332
rect 21980 45444 22036 45454
rect 19740 44994 19796 45006
rect 19740 44942 19742 44994
rect 19794 44942 19796 44994
rect 19740 44660 19796 44942
rect 19740 44594 19796 44604
rect 19852 44884 19908 44894
rect 19404 44436 19460 44446
rect 19292 44434 19460 44436
rect 19292 44382 19406 44434
rect 19458 44382 19460 44434
rect 19292 44380 19460 44382
rect 18396 44212 18452 44222
rect 18396 44118 18452 44156
rect 18732 43764 18788 43774
rect 19292 43764 19348 44380
rect 19404 44370 19460 44380
rect 19852 44322 19908 44828
rect 19852 44270 19854 44322
rect 19906 44270 19908 44322
rect 19852 44258 19908 44270
rect 20076 44322 20132 45276
rect 20076 44270 20078 44322
rect 20130 44270 20132 44322
rect 20076 44258 20132 44270
rect 21868 45108 21924 45118
rect 19516 44100 19572 44110
rect 19964 44100 20020 44110
rect 19516 44006 19572 44044
rect 19628 44098 20020 44100
rect 19628 44046 19966 44098
rect 20018 44046 20020 44098
rect 19628 44044 20020 44046
rect 18732 43650 18788 43708
rect 18732 43598 18734 43650
rect 18786 43598 18788 43650
rect 18732 43586 18788 43598
rect 19180 43708 19292 43764
rect 19628 43764 19684 44044
rect 19964 44034 20020 44044
rect 20300 44100 20356 44110
rect 21868 44100 21924 45052
rect 21980 44324 22036 45388
rect 22652 45106 22708 45500
rect 22652 45054 22654 45106
rect 22706 45054 22708 45106
rect 22652 45042 22708 45054
rect 22092 44548 22148 44558
rect 22092 44546 22708 44548
rect 22092 44494 22094 44546
rect 22146 44494 22708 44546
rect 22092 44492 22708 44494
rect 22092 44482 22148 44492
rect 22204 44324 22260 44334
rect 21980 44322 22260 44324
rect 21980 44270 22206 44322
rect 22258 44270 22260 44322
rect 21980 44268 22260 44270
rect 22204 44258 22260 44268
rect 22540 44212 22596 44222
rect 22540 44118 22596 44156
rect 22092 44100 22148 44110
rect 21868 44044 22092 44100
rect 20300 44006 20356 44044
rect 22092 44006 22148 44044
rect 19836 43932 20100 43942
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 19836 43866 20100 43876
rect 19628 43708 20132 43764
rect 18284 43486 18286 43538
rect 18338 43486 18340 43538
rect 18284 43474 18340 43486
rect 18956 43540 19012 43550
rect 18956 43446 19012 43484
rect 18508 43428 18564 43438
rect 18508 43334 18564 43372
rect 18060 41346 18116 41356
rect 17052 41246 17054 41298
rect 17106 41246 17108 41298
rect 17052 41234 17108 41246
rect 19180 41298 19236 43708
rect 19292 43698 19348 43708
rect 20076 43650 20132 43708
rect 20076 43598 20078 43650
rect 20130 43598 20132 43650
rect 20076 43586 20132 43598
rect 20188 43762 20244 43774
rect 20188 43710 20190 43762
rect 20242 43710 20244 43762
rect 20188 43708 20244 43710
rect 21420 43764 21476 43774
rect 20188 43652 20356 43708
rect 21420 43670 21476 43708
rect 19852 43428 19908 43438
rect 20188 43428 20244 43652
rect 19852 43426 20244 43428
rect 19852 43374 19854 43426
rect 19906 43374 20244 43426
rect 19852 43372 20244 43374
rect 19852 43362 19908 43372
rect 19836 42364 20100 42374
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 19836 42298 20100 42308
rect 19180 41246 19182 41298
rect 19234 41246 19236 41298
rect 18620 40404 18676 40414
rect 18620 40310 18676 40348
rect 19068 40404 19124 40414
rect 19068 40310 19124 40348
rect 17388 39730 17444 39742
rect 17388 39678 17390 39730
rect 17442 39678 17444 39730
rect 17052 39620 17108 39630
rect 16940 39618 17108 39620
rect 16940 39566 17054 39618
rect 17106 39566 17108 39618
rect 16940 39564 17108 39566
rect 16380 38782 16382 38834
rect 16434 38782 16436 38834
rect 16380 38770 16436 38782
rect 16604 38836 16660 38846
rect 16604 38742 16660 38780
rect 15708 38612 16660 38668
rect 15932 38052 15988 38062
rect 15932 37378 15988 37996
rect 15932 37326 15934 37378
rect 15986 37326 15988 37378
rect 15932 37314 15988 37326
rect 15260 37214 15262 37266
rect 15314 37214 15316 37266
rect 15260 37202 15316 37214
rect 15820 37266 15876 37278
rect 16492 37268 16548 37278
rect 15820 37214 15822 37266
rect 15874 37214 15876 37266
rect 15820 37156 15876 37214
rect 16044 37266 16548 37268
rect 16044 37214 16494 37266
rect 16546 37214 16548 37266
rect 16044 37212 16548 37214
rect 16044 37156 16100 37212
rect 16492 37202 16548 37212
rect 15708 37100 16100 37156
rect 15148 36430 15150 36482
rect 15202 36430 15204 36482
rect 15148 36418 15204 36430
rect 15484 36482 15540 36494
rect 15484 36430 15486 36482
rect 15538 36430 15540 36482
rect 15484 36372 15540 36430
rect 15484 36306 15540 36316
rect 15596 36370 15652 36382
rect 15596 36318 15598 36370
rect 15650 36318 15652 36370
rect 11676 35924 11732 35934
rect 11004 35252 11172 35308
rect 9548 34916 9604 34926
rect 9548 34802 9604 34860
rect 9548 34750 9550 34802
rect 9602 34750 9604 34802
rect 9548 34738 9604 34750
rect 9884 34804 9940 34814
rect 9884 34802 10052 34804
rect 9884 34750 9886 34802
rect 9938 34750 10052 34802
rect 9884 34748 10052 34750
rect 9884 34738 9940 34748
rect 9548 33458 9604 33470
rect 9548 33406 9550 33458
rect 9602 33406 9604 33458
rect 9436 33124 9492 33134
rect 9436 33030 9492 33068
rect 9548 32674 9604 33406
rect 9884 33236 9940 33246
rect 9884 32786 9940 33180
rect 9884 32734 9886 32786
rect 9938 32734 9940 32786
rect 9884 32722 9940 32734
rect 9548 32622 9550 32674
rect 9602 32622 9604 32674
rect 9548 32610 9604 32622
rect 9660 32674 9716 32686
rect 9660 32622 9662 32674
rect 9714 32622 9716 32674
rect 9100 32172 9380 32228
rect 9100 31780 9156 32172
rect 9660 32116 9716 32622
rect 9100 31686 9156 31724
rect 9324 32060 9716 32116
rect 9324 31778 9380 32060
rect 9996 31892 10052 34748
rect 10556 34132 10612 34142
rect 10556 34038 10612 34076
rect 11116 34132 11172 35252
rect 11116 34066 11172 34076
rect 11228 34018 11284 34030
rect 11228 33966 11230 34018
rect 11282 33966 11284 34018
rect 11228 33460 11284 33966
rect 11676 33460 11732 35868
rect 14364 34916 14420 34926
rect 14364 34822 14420 34860
rect 14812 34916 14868 34926
rect 14812 34822 14868 34860
rect 15036 34804 15092 34814
rect 14924 34802 15092 34804
rect 14924 34750 15038 34802
rect 15090 34750 15092 34802
rect 14924 34748 15092 34750
rect 13804 34132 13860 34142
rect 13804 34038 13860 34076
rect 10444 33404 10948 33460
rect 10444 33346 10500 33404
rect 10444 33294 10446 33346
rect 10498 33294 10500 33346
rect 10444 33282 10500 33294
rect 10892 33346 10948 33404
rect 10892 33294 10894 33346
rect 10946 33294 10948 33346
rect 10892 33282 10948 33294
rect 11004 33404 11284 33460
rect 11340 33458 11732 33460
rect 11340 33406 11678 33458
rect 11730 33406 11732 33458
rect 11340 33404 11732 33406
rect 9324 31726 9326 31778
rect 9378 31726 9380 31778
rect 9212 31554 9268 31566
rect 9212 31502 9214 31554
rect 9266 31502 9268 31554
rect 9212 31108 9268 31502
rect 9324 31556 9380 31726
rect 9324 31490 9380 31500
rect 9436 31890 10052 31892
rect 9436 31838 9998 31890
rect 10050 31838 10052 31890
rect 9436 31836 10052 31838
rect 9212 31042 9268 31052
rect 9436 30434 9492 31836
rect 9996 31826 10052 31836
rect 10108 33234 10164 33246
rect 10108 33182 10110 33234
rect 10162 33182 10164 33234
rect 9772 31554 9828 31566
rect 9772 31502 9774 31554
rect 9826 31502 9828 31554
rect 9660 30996 9716 31006
rect 9772 30996 9828 31502
rect 9884 31556 9940 31566
rect 9884 31462 9940 31500
rect 10108 31108 10164 33182
rect 10668 33236 10724 33246
rect 10668 33142 10724 33180
rect 10220 33124 10276 33134
rect 10220 32004 10276 33068
rect 10892 33124 10948 33134
rect 11004 33124 11060 33404
rect 11228 33236 11284 33246
rect 11340 33236 11396 33404
rect 11676 33394 11732 33404
rect 13356 34018 13412 34030
rect 13356 33966 13358 34018
rect 13410 33966 13412 34018
rect 11228 33234 11396 33236
rect 11228 33182 11230 33234
rect 11282 33182 11396 33234
rect 11228 33180 11396 33182
rect 11228 33170 11284 33180
rect 10892 33122 11060 33124
rect 10892 33070 10894 33122
rect 10946 33070 11060 33122
rect 10892 33068 11060 33070
rect 10892 33058 10948 33068
rect 13020 32452 13076 32462
rect 13020 32358 13076 32396
rect 10556 32004 10612 32014
rect 10220 31948 10556 32004
rect 10556 31666 10612 31948
rect 13356 32004 13412 33966
rect 14700 33346 14756 33358
rect 14700 33294 14702 33346
rect 14754 33294 14756 33346
rect 13692 32562 13748 32574
rect 13692 32510 13694 32562
rect 13746 32510 13748 32562
rect 13692 32452 13748 32510
rect 13692 32386 13748 32396
rect 14252 32562 14308 32574
rect 14252 32510 14254 32562
rect 14306 32510 14308 32562
rect 11116 31892 11172 31902
rect 10556 31614 10558 31666
rect 10610 31614 10612 31666
rect 10556 31602 10612 31614
rect 10668 31666 10724 31678
rect 10668 31614 10670 31666
rect 10722 31614 10724 31666
rect 10108 31042 10164 31052
rect 10332 31554 10388 31566
rect 10332 31502 10334 31554
rect 10386 31502 10388 31554
rect 9996 30996 10052 31006
rect 9660 30994 9828 30996
rect 9660 30942 9662 30994
rect 9714 30942 9828 30994
rect 9660 30940 9828 30942
rect 9884 30994 10052 30996
rect 9884 30942 9998 30994
rect 10050 30942 10052 30994
rect 9884 30940 10052 30942
rect 9660 30930 9716 30940
rect 9548 30882 9604 30894
rect 9548 30830 9550 30882
rect 9602 30830 9604 30882
rect 9548 30772 9604 30830
rect 9548 30716 9716 30772
rect 9436 30382 9438 30434
rect 9490 30382 9492 30434
rect 9436 30212 9492 30382
rect 9548 30436 9604 30446
rect 9548 30342 9604 30380
rect 9660 30324 9716 30716
rect 9884 30434 9940 30940
rect 9996 30930 10052 30940
rect 10220 30994 10276 31006
rect 10220 30942 10222 30994
rect 10274 30942 10276 30994
rect 9884 30382 9886 30434
rect 9938 30382 9940 30434
rect 9884 30370 9940 30382
rect 9772 30324 9828 30334
rect 9660 30268 9772 30324
rect 9772 30230 9828 30268
rect 10220 30324 10276 30942
rect 10220 30258 10276 30268
rect 9436 30156 9716 30212
rect 9660 28644 9716 30156
rect 10108 29988 10164 29998
rect 10108 29314 10164 29932
rect 10108 29262 10110 29314
rect 10162 29262 10164 29314
rect 10108 29250 10164 29262
rect 10220 28868 10276 28878
rect 10332 28868 10388 31502
rect 10556 31108 10612 31118
rect 10556 31014 10612 31052
rect 10444 30882 10500 30894
rect 10444 30830 10446 30882
rect 10498 30830 10500 30882
rect 10444 29652 10500 30830
rect 10668 30324 10724 31614
rect 10668 30258 10724 30268
rect 11116 30996 11172 31836
rect 11228 30996 11284 31006
rect 11116 30994 11284 30996
rect 11116 30942 11230 30994
rect 11282 30942 11284 30994
rect 11116 30940 11284 30942
rect 11116 30322 11172 30940
rect 11228 30930 11284 30940
rect 12012 30884 12068 30894
rect 11116 30270 11118 30322
rect 11170 30270 11172 30322
rect 11116 30258 11172 30270
rect 11452 30882 12068 30884
rect 11452 30830 12014 30882
rect 12066 30830 12068 30882
rect 11452 30828 12068 30830
rect 10444 29596 11172 29652
rect 10220 28866 10388 28868
rect 10220 28814 10222 28866
rect 10274 28814 10388 28866
rect 10220 28812 10388 28814
rect 10220 28802 10276 28812
rect 9884 28644 9940 28654
rect 9660 28642 10052 28644
rect 9660 28590 9886 28642
rect 9938 28590 10052 28642
rect 9660 28588 10052 28590
rect 9884 28578 9940 28588
rect 8988 28354 9044 28364
rect 8988 27860 9044 27870
rect 9660 27860 9716 27870
rect 8988 27858 9716 27860
rect 8988 27806 8990 27858
rect 9042 27806 9662 27858
rect 9714 27806 9716 27858
rect 8988 27804 9716 27806
rect 9996 27860 10052 28588
rect 10108 28420 10164 28430
rect 10108 28418 10276 28420
rect 10108 28366 10110 28418
rect 10162 28366 10276 28418
rect 10108 28364 10276 28366
rect 10108 28354 10164 28364
rect 10108 27860 10164 27870
rect 9996 27858 10164 27860
rect 9996 27806 10110 27858
rect 10162 27806 10164 27858
rect 9996 27804 10164 27806
rect 8988 27794 9044 27804
rect 9660 27794 9716 27804
rect 10108 27794 10164 27804
rect 8876 27746 8932 27758
rect 8876 27694 8878 27746
rect 8930 27694 8932 27746
rect 8876 27636 8932 27694
rect 8876 27580 9044 27636
rect 8988 27076 9044 27580
rect 8988 27010 9044 27020
rect 9548 27634 9604 27646
rect 9548 27582 9550 27634
rect 9602 27582 9604 27634
rect 8540 25666 8596 25676
rect 8652 26852 8820 26908
rect 8876 26964 8932 26974
rect 8428 25218 8484 25228
rect 8540 25506 8596 25518
rect 8540 25454 8542 25506
rect 8594 25454 8596 25506
rect 8540 23940 8596 25454
rect 8652 25396 8708 26852
rect 8764 26404 8820 26414
rect 8876 26404 8932 26908
rect 8764 26402 8932 26404
rect 8764 26350 8766 26402
rect 8818 26350 8932 26402
rect 8764 26348 8932 26350
rect 8764 25732 8820 26348
rect 9548 26292 9604 27582
rect 9772 27076 9828 27086
rect 9772 26962 9828 27020
rect 10220 27076 10276 28364
rect 10332 27858 10388 28812
rect 11116 28866 11172 29596
rect 11116 28814 11118 28866
rect 11170 28814 11172 28866
rect 11116 28802 11172 28814
rect 11452 28866 11508 30828
rect 12012 30818 12068 30828
rect 12796 30210 12852 30222
rect 12796 30158 12798 30210
rect 12850 30158 12852 30210
rect 12796 29652 12852 30158
rect 13356 30212 13412 31948
rect 14252 31892 14308 32510
rect 14364 32564 14420 32574
rect 14364 32470 14420 32508
rect 14588 31892 14644 31902
rect 14252 31836 14588 31892
rect 14588 31798 14644 31836
rect 13580 31556 13636 31566
rect 13356 30146 13412 30156
rect 13468 30324 13524 30334
rect 13468 30098 13524 30268
rect 13468 30046 13470 30098
rect 13522 30046 13524 30098
rect 13468 30034 13524 30046
rect 13020 29652 13076 29662
rect 13468 29652 13524 29662
rect 13580 29652 13636 31500
rect 14140 30996 14196 31006
rect 14140 30884 14196 30940
rect 13804 30882 14196 30884
rect 13804 30830 14142 30882
rect 14194 30830 14196 30882
rect 13804 30828 14196 30830
rect 13804 30210 13860 30828
rect 14140 30818 14196 30828
rect 13804 30158 13806 30210
rect 13858 30158 13860 30210
rect 13804 30146 13860 30158
rect 12348 29650 13636 29652
rect 12348 29598 13022 29650
rect 13074 29598 13470 29650
rect 13522 29598 13636 29650
rect 12348 29596 13636 29598
rect 12348 29426 12404 29596
rect 13020 29586 13076 29596
rect 13468 29586 13524 29596
rect 12348 29374 12350 29426
rect 12402 29374 12404 29426
rect 12348 29362 12404 29374
rect 11452 28814 11454 28866
rect 11506 28814 11508 28866
rect 11452 28802 11508 28814
rect 11340 28644 11396 28654
rect 11340 28530 11396 28588
rect 11900 28644 11956 28654
rect 11900 28550 11956 28588
rect 11340 28478 11342 28530
rect 11394 28478 11396 28530
rect 11340 28466 11396 28478
rect 10444 28082 10500 28094
rect 10444 28030 10446 28082
rect 10498 28030 10500 28082
rect 10444 27972 10500 28030
rect 11564 28084 11620 28094
rect 11564 27990 11620 28028
rect 12684 28084 12740 28094
rect 10780 27972 10836 27982
rect 10444 27970 10836 27972
rect 10444 27918 10782 27970
rect 10834 27918 10836 27970
rect 10444 27916 10836 27918
rect 10332 27806 10334 27858
rect 10386 27806 10388 27858
rect 10332 27794 10388 27806
rect 10444 27076 10500 27086
rect 10220 27074 10500 27076
rect 10220 27022 10222 27074
rect 10274 27022 10446 27074
rect 10498 27022 10500 27074
rect 10220 27020 10500 27022
rect 10220 27010 10276 27020
rect 10444 27010 10500 27020
rect 9772 26910 9774 26962
rect 9826 26910 9828 26962
rect 9772 26898 9828 26910
rect 9996 26964 10052 27002
rect 9996 26898 10052 26908
rect 9548 26226 9604 26236
rect 9660 26850 9716 26862
rect 9660 26798 9662 26850
rect 9714 26798 9716 26850
rect 8764 25676 9380 25732
rect 8652 25330 8708 25340
rect 8764 24052 8820 24062
rect 8316 23884 8484 23940
rect 8204 23828 8260 23884
rect 8092 23826 8260 23828
rect 8092 23774 8206 23826
rect 8258 23774 8260 23826
rect 8092 23772 8260 23774
rect 7980 23716 8036 23726
rect 7868 23714 8036 23716
rect 7868 23662 7982 23714
rect 8034 23662 8036 23714
rect 7868 23660 8036 23662
rect 7868 23380 7924 23660
rect 7980 23650 8036 23660
rect 7644 23324 7924 23380
rect 7644 23268 7700 23324
rect 7644 23174 7700 23212
rect 7868 23156 7924 23166
rect 8092 23156 8148 23772
rect 8204 23762 8260 23772
rect 8316 23716 8372 23726
rect 8316 23622 8372 23660
rect 8428 23492 8484 23884
rect 8540 23874 8596 23884
rect 8652 24050 8820 24052
rect 8652 23998 8766 24050
rect 8818 23998 8820 24050
rect 8652 23996 8820 23998
rect 7868 23154 8148 23156
rect 7868 23102 7870 23154
rect 7922 23102 8148 23154
rect 7868 23100 8148 23102
rect 8316 23436 8484 23492
rect 7868 23090 7924 23100
rect 7420 23044 7476 23054
rect 7420 22950 7476 22988
rect 8092 21812 8148 21822
rect 8092 21718 8148 21756
rect 8316 21810 8372 23436
rect 8428 23154 8484 23166
rect 8428 23102 8430 23154
rect 8482 23102 8484 23154
rect 8428 23044 8484 23102
rect 8652 23154 8708 23996
rect 8764 23986 8820 23996
rect 8876 23940 8932 23950
rect 8876 23846 8932 23884
rect 8764 23828 8820 23838
rect 8764 23734 8820 23772
rect 9324 23826 9380 25676
rect 9436 25506 9492 25518
rect 9436 25454 9438 25506
rect 9490 25454 9492 25506
rect 9436 25284 9492 25454
rect 9660 25508 9716 26798
rect 9660 25442 9716 25452
rect 10556 25506 10612 27916
rect 10780 27906 10836 27916
rect 11004 27972 11060 27982
rect 11004 27878 11060 27916
rect 12684 27970 12740 28028
rect 12684 27918 12686 27970
rect 12738 27918 12740 27970
rect 12684 27906 12740 27918
rect 11564 27858 11620 27870
rect 11900 27860 11956 27870
rect 11564 27806 11566 27858
rect 11618 27806 11620 27858
rect 11228 27636 11284 27646
rect 10668 27634 11284 27636
rect 10668 27582 11230 27634
rect 11282 27582 11284 27634
rect 10668 27580 11284 27582
rect 10668 27186 10724 27580
rect 11228 27570 11284 27580
rect 10668 27134 10670 27186
rect 10722 27134 10724 27186
rect 10668 27122 10724 27134
rect 11564 27188 11620 27806
rect 11564 27122 11620 27132
rect 11676 27858 11956 27860
rect 11676 27806 11902 27858
rect 11954 27806 11956 27858
rect 11676 27804 11956 27806
rect 10780 27074 10836 27086
rect 10780 27022 10782 27074
rect 10834 27022 10836 27074
rect 10780 26964 10836 27022
rect 11116 27076 11172 27086
rect 11116 26982 11172 27020
rect 10780 26898 10836 26908
rect 11676 26964 11732 27804
rect 11900 27794 11956 27804
rect 14700 27748 14756 33294
rect 14812 32564 14868 32574
rect 14924 32564 14980 34748
rect 15036 34738 15092 34748
rect 15484 34692 15540 34702
rect 15484 34598 15540 34636
rect 15596 34356 15652 36318
rect 15148 34300 15652 34356
rect 15036 33348 15092 33358
rect 15036 33012 15092 33292
rect 15036 32946 15092 32956
rect 15036 32564 15092 32574
rect 14924 32562 15092 32564
rect 14924 32510 15038 32562
rect 15090 32510 15092 32562
rect 14924 32508 15092 32510
rect 15148 32564 15204 34300
rect 15484 34132 15540 34142
rect 15708 34132 15764 37100
rect 16268 37044 16324 37054
rect 16044 36372 16100 36382
rect 16044 36278 16100 36316
rect 16268 35698 16324 36988
rect 16604 35812 16660 38612
rect 16268 35646 16270 35698
rect 16322 35646 16324 35698
rect 16268 35634 16324 35646
rect 16492 35756 16660 35812
rect 15484 34130 15764 34132
rect 15484 34078 15486 34130
rect 15538 34078 15764 34130
rect 15484 34076 15764 34078
rect 15820 35586 15876 35598
rect 15820 35534 15822 35586
rect 15874 35534 15876 35586
rect 15484 33572 15540 34076
rect 15484 33506 15540 33516
rect 15260 33236 15316 33246
rect 15260 33234 15540 33236
rect 15260 33182 15262 33234
rect 15314 33182 15540 33234
rect 15260 33180 15540 33182
rect 15260 33170 15316 33180
rect 15372 33012 15428 33022
rect 15260 32564 15316 32574
rect 15148 32562 15316 32564
rect 15148 32510 15262 32562
rect 15314 32510 15316 32562
rect 15148 32508 15316 32510
rect 14812 32470 14868 32508
rect 15036 32498 15092 32508
rect 15260 32498 15316 32508
rect 15372 32340 15428 32956
rect 15484 32562 15540 33180
rect 15820 32900 15876 35534
rect 15820 32844 16324 32900
rect 16156 32676 16212 32686
rect 16156 32582 16212 32620
rect 15484 32510 15486 32562
rect 15538 32510 15540 32562
rect 15484 32498 15540 32510
rect 15596 32564 15652 32574
rect 16044 32564 16100 32574
rect 15596 32562 16100 32564
rect 15596 32510 15598 32562
rect 15650 32510 16046 32562
rect 16098 32510 16100 32562
rect 15596 32508 16100 32510
rect 15596 32498 15652 32508
rect 16044 32498 16100 32508
rect 15148 32284 15428 32340
rect 16268 32340 16324 32844
rect 16380 32562 16436 32574
rect 16380 32510 16382 32562
rect 16434 32510 16436 32562
rect 16380 32452 16436 32510
rect 16492 32564 16548 35756
rect 16604 35588 16660 35598
rect 16604 35494 16660 35532
rect 16604 34692 16660 34702
rect 16604 32788 16660 34636
rect 16716 33458 16772 39564
rect 17052 39554 17108 39564
rect 16828 38722 16884 38734
rect 16828 38670 16830 38722
rect 16882 38670 16884 38722
rect 16828 38388 16884 38670
rect 16828 38322 16884 38332
rect 17388 38722 17444 39678
rect 18956 39620 19012 39630
rect 19180 39620 19236 41246
rect 19516 41636 19572 41646
rect 18956 39618 19236 39620
rect 18956 39566 18958 39618
rect 19010 39566 19236 39618
rect 18956 39564 19236 39566
rect 19292 39618 19348 39630
rect 19292 39566 19294 39618
rect 19346 39566 19348 39618
rect 18956 39554 19012 39564
rect 17724 39506 17780 39518
rect 17724 39454 17726 39506
rect 17778 39454 17780 39506
rect 17388 38670 17390 38722
rect 17442 38670 17444 38722
rect 16716 33406 16718 33458
rect 16770 33406 16772 33458
rect 16716 33394 16772 33406
rect 16604 32722 16660 32732
rect 16492 32508 16660 32564
rect 16380 32396 16548 32452
rect 16268 32284 16436 32340
rect 14812 29652 14868 29662
rect 14812 29426 14868 29596
rect 14812 29374 14814 29426
rect 14866 29374 14868 29426
rect 14812 29362 14868 29374
rect 14812 27748 14868 27758
rect 14700 27746 14868 27748
rect 14700 27694 14814 27746
rect 14866 27694 14868 27746
rect 14700 27692 14868 27694
rect 11788 27188 11844 27198
rect 11788 27094 11844 27132
rect 14700 27076 14756 27692
rect 14812 27682 14868 27692
rect 14700 27010 14756 27020
rect 10556 25454 10558 25506
rect 10610 25454 10612 25506
rect 10556 25442 10612 25454
rect 10780 25506 10836 25518
rect 10780 25454 10782 25506
rect 10834 25454 10836 25506
rect 9884 25284 9940 25294
rect 9436 25282 10052 25284
rect 9436 25230 9886 25282
rect 9938 25230 10052 25282
rect 9436 25228 10052 25230
rect 9884 25218 9940 25228
rect 9324 23774 9326 23826
rect 9378 23774 9380 23826
rect 8652 23102 8654 23154
rect 8706 23102 8708 23154
rect 8652 23090 8708 23102
rect 9100 23716 9156 23726
rect 8428 22978 8484 22988
rect 8988 23044 9044 23054
rect 8988 22950 9044 22988
rect 8876 22932 8932 22942
rect 8316 21758 8318 21810
rect 8370 21758 8372 21810
rect 8316 21746 8372 21758
rect 8652 21812 8708 21822
rect 7980 21586 8036 21598
rect 7980 21534 7982 21586
rect 8034 21534 8036 21586
rect 7532 21028 7588 21038
rect 7308 21026 7588 21028
rect 7308 20974 7534 21026
rect 7586 20974 7588 21026
rect 7308 20972 7588 20974
rect 7532 20962 7588 20972
rect 7868 20692 7924 20702
rect 7980 20692 8036 21534
rect 7868 20690 8036 20692
rect 7868 20638 7870 20690
rect 7922 20638 8036 20690
rect 7868 20636 8036 20638
rect 8652 21474 8708 21756
rect 8652 21422 8654 21474
rect 8706 21422 8708 21474
rect 7644 20578 7700 20590
rect 7644 20526 7646 20578
rect 7698 20526 7700 20578
rect 6860 20078 6862 20130
rect 6914 20078 6916 20130
rect 6860 20066 6916 20078
rect 7084 20132 7140 20142
rect 6412 20018 6468 20030
rect 7084 20020 7140 20076
rect 6412 19966 6414 20018
rect 6466 19966 6468 20018
rect 4956 19908 5012 19918
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 4956 19458 5012 19852
rect 6412 19908 6468 19966
rect 6412 19842 6468 19852
rect 6972 20018 7140 20020
rect 6972 19966 7086 20018
rect 7138 19966 7140 20018
rect 6972 19964 7140 19966
rect 6972 19460 7028 19964
rect 7084 19954 7140 19964
rect 7308 20020 7364 20030
rect 7644 20020 7700 20526
rect 7868 20244 7924 20636
rect 8652 20468 8708 21422
rect 8652 20402 8708 20412
rect 8764 20692 8820 20702
rect 7868 20188 8260 20244
rect 7308 20018 7588 20020
rect 7308 19966 7310 20018
rect 7362 19966 7588 20018
rect 7308 19964 7588 19966
rect 7644 19964 8148 20020
rect 7308 19954 7364 19964
rect 4956 19406 4958 19458
rect 5010 19406 5012 19458
rect 4956 19394 5012 19406
rect 6860 19404 7028 19460
rect 7084 19796 7140 19806
rect 7084 19458 7140 19740
rect 7084 19406 7086 19458
rect 7138 19406 7140 19458
rect 5628 19234 5684 19246
rect 5628 19182 5630 19234
rect 5682 19182 5684 19234
rect 5068 19122 5124 19134
rect 5068 19070 5070 19122
rect 5122 19070 5124 19122
rect 4956 19012 5012 19022
rect 1820 18450 1876 18462
rect 1820 18398 1822 18450
rect 1874 18398 1876 18450
rect 1820 16884 1876 18398
rect 2492 18452 2548 18462
rect 2492 18358 2548 18396
rect 4620 18340 4676 18350
rect 4956 18340 5012 18956
rect 5068 18788 5124 19070
rect 5628 19012 5684 19182
rect 5628 18946 5684 18956
rect 5852 19234 5908 19246
rect 5852 19182 5854 19234
rect 5906 19182 5908 19234
rect 5852 18788 5908 19182
rect 6524 19122 6580 19134
rect 6524 19070 6526 19122
rect 6578 19070 6580 19122
rect 6188 19012 6244 19022
rect 6188 18918 6244 18956
rect 5068 18732 5908 18788
rect 5516 18450 5572 18462
rect 5516 18398 5518 18450
rect 5570 18398 5572 18450
rect 5068 18340 5124 18350
rect 4956 18338 5124 18340
rect 4956 18286 5070 18338
rect 5122 18286 5124 18338
rect 4956 18284 5124 18286
rect 4620 18246 4676 18284
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 5068 17892 5124 18284
rect 4620 17836 5124 17892
rect 5516 18340 5572 18398
rect 4620 17106 4676 17836
rect 5516 17556 5572 18284
rect 5516 17490 5572 17500
rect 4620 17054 4622 17106
rect 4674 17054 4676 17106
rect 4620 17042 4676 17054
rect 4844 17442 4900 17454
rect 4844 17390 4846 17442
rect 4898 17390 4900 17442
rect 1820 16098 1876 16828
rect 4732 16994 4788 17006
rect 4732 16942 4734 16994
rect 4786 16942 4788 16994
rect 4508 16660 4564 16670
rect 4284 16658 4564 16660
rect 4284 16606 4510 16658
rect 4562 16606 4564 16658
rect 4284 16604 4564 16606
rect 4732 16660 4788 16942
rect 4844 16884 4900 17390
rect 5068 16884 5124 16894
rect 4844 16828 5068 16884
rect 4732 16604 5012 16660
rect 4284 16324 4340 16604
rect 4508 16594 4564 16604
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 4284 16268 4676 16324
rect 1820 16046 1822 16098
rect 1874 16046 1876 16098
rect 1820 16034 1876 16046
rect 4620 16210 4676 16268
rect 4620 16158 4622 16210
rect 4674 16158 4676 16210
rect 2492 15988 2548 15998
rect 2268 15986 2548 15988
rect 2268 15934 2494 15986
rect 2546 15934 2548 15986
rect 2268 15932 2548 15934
rect 2268 15538 2324 15932
rect 2492 15922 2548 15932
rect 2268 15486 2270 15538
rect 2322 15486 2324 15538
rect 2268 15474 2324 15486
rect 4620 15538 4676 16158
rect 4956 16100 5012 16604
rect 5068 16210 5124 16828
rect 5068 16158 5070 16210
rect 5122 16158 5124 16210
rect 5068 16146 5124 16158
rect 4620 15486 4622 15538
rect 4674 15486 4676 15538
rect 4620 15474 4676 15486
rect 4844 16044 5012 16100
rect 2604 15316 2660 15326
rect 2604 15222 2660 15260
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 4844 13972 4900 16044
rect 5852 15988 5908 18732
rect 6412 18562 6468 18574
rect 6412 18510 6414 18562
rect 6466 18510 6468 18562
rect 5964 18452 6020 18462
rect 6300 18452 6356 18462
rect 5964 18450 6356 18452
rect 5964 18398 5966 18450
rect 6018 18398 6302 18450
rect 6354 18398 6356 18450
rect 5964 18396 6356 18398
rect 5964 18386 6020 18396
rect 6300 18386 6356 18396
rect 6412 17780 6468 18510
rect 6412 17714 6468 17724
rect 6524 17778 6580 19070
rect 6748 19122 6804 19134
rect 6748 19070 6750 19122
rect 6802 19070 6804 19122
rect 6636 19010 6692 19022
rect 6636 18958 6638 19010
rect 6690 18958 6692 19010
rect 6636 18900 6692 18958
rect 6636 18834 6692 18844
rect 6748 18676 6804 19070
rect 6860 19012 6916 19404
rect 7084 19394 7140 19406
rect 7084 19234 7140 19246
rect 7084 19182 7086 19234
rect 7138 19182 7140 19234
rect 7084 19124 7140 19182
rect 7532 19124 7588 19964
rect 8092 19906 8148 19964
rect 8092 19854 8094 19906
rect 8146 19854 8148 19906
rect 7644 19796 7700 19806
rect 7700 19740 7812 19796
rect 7644 19730 7700 19740
rect 7644 19124 7700 19134
rect 7084 19058 7140 19068
rect 7196 19122 7700 19124
rect 7196 19070 7646 19122
rect 7698 19070 7700 19122
rect 7196 19068 7700 19070
rect 6860 18956 7028 19012
rect 6636 18620 6804 18676
rect 6636 18450 6692 18620
rect 6636 18398 6638 18450
rect 6690 18398 6692 18450
rect 6636 18386 6692 18398
rect 6972 18228 7028 18956
rect 6524 17726 6526 17778
rect 6578 17726 6580 17778
rect 6524 17714 6580 17726
rect 6636 18172 7028 18228
rect 6300 17556 6356 17566
rect 5964 16098 6020 16110
rect 5964 16046 5966 16098
rect 6018 16046 6020 16098
rect 5964 15988 6020 16046
rect 6188 16100 6244 16110
rect 6188 16006 6244 16044
rect 5740 15932 6020 15988
rect 4956 15428 5012 15438
rect 4956 15334 5012 15372
rect 5740 15148 5796 15932
rect 5068 15092 5796 15148
rect 4844 13916 5012 13972
rect 2492 13636 2548 13646
rect 2492 13074 2548 13580
rect 4844 13522 4900 13534
rect 4844 13470 4846 13522
rect 4898 13470 4900 13522
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4844 13300 4900 13470
rect 4844 13234 4900 13244
rect 2492 13022 2494 13074
rect 2546 13022 2548 13074
rect 2492 13010 2548 13022
rect 4620 13076 4676 13086
rect 4956 13076 5012 13916
rect 5068 13634 5124 15092
rect 6188 14308 6244 14318
rect 5068 13582 5070 13634
rect 5122 13582 5124 13634
rect 5068 13570 5124 13582
rect 5180 13746 5236 13758
rect 5180 13694 5182 13746
rect 5234 13694 5236 13746
rect 4620 13074 4956 13076
rect 4620 13022 4622 13074
rect 4674 13022 4956 13074
rect 4620 13020 4956 13022
rect 4620 13010 4676 13020
rect 4956 12982 5012 13020
rect 1820 12962 1876 12974
rect 1820 12910 1822 12962
rect 1874 12910 1876 12962
rect 1820 12068 1876 12910
rect 5068 12964 5124 12974
rect 5068 12870 5124 12908
rect 4956 12852 5012 12862
rect 4956 12740 5012 12796
rect 5180 12740 5236 13694
rect 5964 13746 6020 13758
rect 5964 13694 5966 13746
rect 6018 13694 6020 13746
rect 5740 13076 5796 13086
rect 5740 12962 5796 13020
rect 5740 12910 5742 12962
rect 5794 12910 5796 12962
rect 5740 12898 5796 12910
rect 5964 12964 6020 13694
rect 6188 13746 6244 14252
rect 6188 13694 6190 13746
rect 6242 13694 6244 13746
rect 6188 13682 6244 13694
rect 6076 13636 6132 13646
rect 6076 13542 6132 13580
rect 6300 13300 6356 17500
rect 6412 17554 6468 17566
rect 6412 17502 6414 17554
rect 6466 17502 6468 17554
rect 6412 16548 6468 17502
rect 6412 16482 6468 16492
rect 6524 17556 6580 17566
rect 6636 17556 6692 18172
rect 7196 18004 7252 19068
rect 7644 19058 7700 19068
rect 7644 18676 7700 18686
rect 7756 18676 7812 19740
rect 7980 19794 8036 19806
rect 7980 19742 7982 19794
rect 8034 19742 8036 19794
rect 7980 19348 8036 19742
rect 7980 19234 8036 19292
rect 7980 19182 7982 19234
rect 8034 19182 8036 19234
rect 7980 19170 8036 19182
rect 7644 18674 7812 18676
rect 7644 18622 7646 18674
rect 7698 18622 7812 18674
rect 7644 18620 7812 18622
rect 7644 18610 7700 18620
rect 8092 18340 8148 19854
rect 8204 19124 8260 20188
rect 8652 20132 8708 20142
rect 8652 20038 8708 20076
rect 8316 20020 8372 20030
rect 8316 19926 8372 19964
rect 8540 19348 8596 19358
rect 8540 19254 8596 19292
rect 8316 19124 8372 19134
rect 8204 19068 8316 19124
rect 8316 19058 8372 19068
rect 6748 17948 7252 18004
rect 7868 18284 8148 18340
rect 6748 17666 6804 17948
rect 6748 17614 6750 17666
rect 6802 17614 6804 17666
rect 6748 17602 6804 17614
rect 6972 17780 7028 17790
rect 6524 17554 6692 17556
rect 6524 17502 6526 17554
rect 6578 17502 6692 17554
rect 6524 17500 6692 17502
rect 6412 16324 6468 16334
rect 6524 16324 6580 17500
rect 6412 16322 6580 16324
rect 6412 16270 6414 16322
rect 6466 16270 6580 16322
rect 6412 16268 6580 16270
rect 6412 16258 6468 16268
rect 6524 16212 6580 16268
rect 6524 16146 6580 16156
rect 6524 15986 6580 15998
rect 6524 15934 6526 15986
rect 6578 15934 6580 15986
rect 6524 14532 6580 15934
rect 6972 14868 7028 17724
rect 7084 16100 7140 17948
rect 7644 17444 7700 17454
rect 7868 17444 7924 18284
rect 7980 17780 8036 17790
rect 7980 17554 8036 17724
rect 7980 17502 7982 17554
rect 8034 17502 8036 17554
rect 7980 17490 8036 17502
rect 7644 17442 7924 17444
rect 7644 17390 7646 17442
rect 7698 17390 7924 17442
rect 7644 17388 7924 17390
rect 7644 17220 7700 17388
rect 7084 16034 7140 16044
rect 7196 17164 7700 17220
rect 7084 15428 7140 15438
rect 7084 15334 7140 15372
rect 7196 15426 7252 17164
rect 7532 16212 7588 16222
rect 7308 16100 7364 16110
rect 7308 16006 7364 16044
rect 7532 16098 7588 16156
rect 7532 16046 7534 16098
rect 7586 16046 7588 16098
rect 7532 16034 7588 16046
rect 7980 16100 8036 16110
rect 7980 16098 8596 16100
rect 7980 16046 7982 16098
rect 8034 16046 8596 16098
rect 7980 16044 8596 16046
rect 7980 16034 8036 16044
rect 7420 15874 7476 15886
rect 7420 15822 7422 15874
rect 7474 15822 7476 15874
rect 7420 15540 7476 15822
rect 7420 15484 8260 15540
rect 7196 15374 7198 15426
rect 7250 15374 7252 15426
rect 7196 15362 7252 15374
rect 8204 15426 8260 15484
rect 8540 15538 8596 16044
rect 8764 15652 8820 20636
rect 8876 19796 8932 22876
rect 9100 21252 9156 23660
rect 9324 23268 9380 23774
rect 9772 25060 9828 25070
rect 9772 23378 9828 25004
rect 9772 23326 9774 23378
rect 9826 23326 9828 23378
rect 9772 23314 9828 23326
rect 9548 23268 9604 23278
rect 9324 23266 9604 23268
rect 9324 23214 9550 23266
rect 9602 23214 9604 23266
rect 9324 23212 9604 23214
rect 9548 23202 9604 23212
rect 9996 23154 10052 25228
rect 10668 24834 10724 24846
rect 10668 24782 10670 24834
rect 10722 24782 10724 24834
rect 10668 24724 10724 24782
rect 10668 24658 10724 24668
rect 9996 23102 9998 23154
rect 10050 23102 10052 23154
rect 9884 23042 9940 23054
rect 9884 22990 9886 23042
rect 9938 22990 9940 23042
rect 9212 22932 9268 22942
rect 9212 22482 9268 22876
rect 9212 22430 9214 22482
rect 9266 22430 9268 22482
rect 9212 22418 9268 22430
rect 9660 21812 9716 21822
rect 9660 21718 9716 21756
rect 9884 21700 9940 22990
rect 9996 21924 10052 23102
rect 10108 24612 10164 24622
rect 10108 22820 10164 24556
rect 10780 24610 10836 25454
rect 10780 24558 10782 24610
rect 10834 24558 10836 24610
rect 10780 24546 10836 24558
rect 11004 25506 11060 25518
rect 11004 25454 11006 25506
rect 11058 25454 11060 25506
rect 11004 25284 11060 25454
rect 11116 25508 11172 25546
rect 11116 25442 11172 25452
rect 11564 25506 11620 25518
rect 11564 25454 11566 25506
rect 11618 25454 11620 25506
rect 10444 24500 10500 24510
rect 10444 24498 10612 24500
rect 10444 24446 10446 24498
rect 10498 24446 10612 24498
rect 10444 24444 10612 24446
rect 10444 24434 10500 24444
rect 10556 23828 10612 24444
rect 10556 23378 10612 23772
rect 10556 23326 10558 23378
rect 10610 23326 10612 23378
rect 10556 23314 10612 23326
rect 10220 23154 10276 23166
rect 10220 23102 10222 23154
rect 10274 23102 10276 23154
rect 10220 23044 10276 23102
rect 10780 23154 10836 23166
rect 10780 23102 10782 23154
rect 10834 23102 10836 23154
rect 10780 23044 10836 23102
rect 10220 22988 10836 23044
rect 10108 22764 10500 22820
rect 9996 21858 10052 21868
rect 9884 21644 10276 21700
rect 9996 21476 10052 21486
rect 10220 21476 10276 21644
rect 10444 21586 10500 22764
rect 10444 21534 10446 21586
rect 10498 21534 10500 21586
rect 10444 21522 10500 21534
rect 10220 21420 10388 21476
rect 9996 21382 10052 21420
rect 10108 21364 10164 21374
rect 10108 21362 10276 21364
rect 10108 21310 10110 21362
rect 10162 21310 10276 21362
rect 10108 21308 10276 21310
rect 10108 21298 10164 21308
rect 9100 21196 10052 21252
rect 9884 21028 9940 21038
rect 9660 20468 9716 20478
rect 9548 20412 9660 20468
rect 8876 19730 8932 19740
rect 8988 20020 9044 20030
rect 8988 19460 9044 19964
rect 8988 19394 9044 19404
rect 9100 19348 9156 19358
rect 8988 19236 9044 19246
rect 9100 19236 9156 19292
rect 8988 19234 9156 19236
rect 8988 19182 8990 19234
rect 9042 19182 9156 19234
rect 8988 19180 9156 19182
rect 8988 19170 9044 19180
rect 8540 15486 8542 15538
rect 8594 15486 8596 15538
rect 8540 15474 8596 15486
rect 8652 15596 8820 15652
rect 8204 15374 8206 15426
rect 8258 15374 8260 15426
rect 8204 15362 8260 15374
rect 8316 15428 8372 15438
rect 7532 15316 7588 15326
rect 7532 15222 7588 15260
rect 7980 15314 8036 15326
rect 7980 15262 7982 15314
rect 8034 15262 8036 15314
rect 7980 15148 8036 15262
rect 8092 15316 8148 15326
rect 8092 15222 8148 15260
rect 7084 15092 7140 15102
rect 7644 15092 8036 15148
rect 7084 15090 7700 15092
rect 7084 15038 7086 15090
rect 7138 15038 7700 15090
rect 7084 15036 7700 15038
rect 7084 15026 7140 15036
rect 6972 14812 7140 14868
rect 7084 14644 7140 14812
rect 7084 14588 7476 14644
rect 6972 14532 7028 14542
rect 6524 14530 7028 14532
rect 6524 14478 6974 14530
rect 7026 14478 7028 14530
rect 6524 14476 7028 14478
rect 6972 14466 7028 14476
rect 7084 14308 7140 14318
rect 7084 14214 7140 14252
rect 7196 14306 7252 14318
rect 7196 14254 7198 14306
rect 7250 14254 7252 14306
rect 6412 13972 6468 13982
rect 6412 13746 6468 13916
rect 6412 13694 6414 13746
rect 6466 13694 6468 13746
rect 6412 13682 6468 13694
rect 6636 13746 6692 13758
rect 6636 13694 6638 13746
rect 6690 13694 6692 13746
rect 6412 13300 6468 13310
rect 6300 13244 6412 13300
rect 6636 13300 6692 13694
rect 6972 13748 7028 13758
rect 6972 13746 7140 13748
rect 6972 13694 6974 13746
rect 7026 13694 7140 13746
rect 6972 13692 7140 13694
rect 6972 13682 7028 13692
rect 7084 13522 7140 13692
rect 7084 13470 7086 13522
rect 7138 13470 7140 13522
rect 7084 13458 7140 13470
rect 7196 13524 7252 14254
rect 7196 13458 7252 13468
rect 7308 13972 7364 13982
rect 7308 13300 7364 13916
rect 7420 13524 7476 14588
rect 7532 14530 7588 15036
rect 7532 14478 7534 14530
rect 7586 14478 7588 14530
rect 7532 14466 7588 14478
rect 8092 14308 8148 14318
rect 8092 13524 8148 14252
rect 7420 13522 8036 13524
rect 7420 13470 7422 13522
rect 7474 13470 8036 13522
rect 7420 13468 8036 13470
rect 7420 13458 7476 13468
rect 6636 13244 6916 13300
rect 6188 13188 6244 13198
rect 6188 13094 6244 13132
rect 6412 13186 6468 13244
rect 6412 13134 6414 13186
rect 6466 13134 6468 13186
rect 6412 13122 6468 13134
rect 6860 13186 6916 13244
rect 6860 13134 6862 13186
rect 6914 13134 6916 13186
rect 6860 13122 6916 13134
rect 6972 13244 7364 13300
rect 5964 12898 6020 12908
rect 6860 12964 6916 12974
rect 6860 12870 6916 12908
rect 5628 12852 5684 12862
rect 5628 12758 5684 12796
rect 4956 12684 5236 12740
rect 5964 12740 6020 12750
rect 6524 12740 6580 12750
rect 1820 10610 1876 12012
rect 4844 12068 4900 12078
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4844 11396 4900 12012
rect 4620 11340 4900 11396
rect 4284 11284 4340 11294
rect 2492 11172 2548 11182
rect 2492 10722 2548 11116
rect 2492 10670 2494 10722
rect 2546 10670 2548 10722
rect 2492 10658 2548 10670
rect 4172 10836 4228 10846
rect 1820 10558 1822 10610
rect 1874 10558 1876 10610
rect 1820 10546 1876 10558
rect 4172 9828 4228 10780
rect 4284 10052 4340 11228
rect 4620 10836 4676 11340
rect 4956 11282 5012 12684
rect 5852 12292 5908 12302
rect 5852 11506 5908 12236
rect 5852 11454 5854 11506
rect 5906 11454 5908 11506
rect 5852 11442 5908 11454
rect 5964 11508 6020 12684
rect 5964 11442 6020 11452
rect 6300 12738 6580 12740
rect 6300 12686 6526 12738
rect 6578 12686 6580 12738
rect 6300 12684 6580 12686
rect 6076 11394 6132 11406
rect 6076 11342 6078 11394
rect 6130 11342 6132 11394
rect 4956 11230 4958 11282
rect 5010 11230 5012 11282
rect 4956 11172 5012 11230
rect 5068 11284 5124 11294
rect 5628 11284 5684 11294
rect 5068 11282 5684 11284
rect 5068 11230 5070 11282
rect 5122 11230 5630 11282
rect 5682 11230 5684 11282
rect 5068 11228 5684 11230
rect 5068 11218 5124 11228
rect 5628 11218 5684 11228
rect 4620 10770 4676 10780
rect 4732 11116 5012 11172
rect 5740 11172 5796 11182
rect 4620 10500 4676 10510
rect 4732 10500 4788 11116
rect 5740 11078 5796 11116
rect 6076 11172 6132 11342
rect 6300 11394 6356 12684
rect 6524 12674 6580 12684
rect 6300 11342 6302 11394
rect 6354 11342 6356 11394
rect 6300 11330 6356 11342
rect 6636 11396 6692 11406
rect 6636 11302 6692 11340
rect 6076 11106 6132 11116
rect 6972 11172 7028 13244
rect 7196 13076 7252 13086
rect 7196 12982 7252 13020
rect 7868 12068 7924 12078
rect 7308 12066 7924 12068
rect 7308 12014 7870 12066
rect 7922 12014 7924 12066
rect 7308 12012 7924 12014
rect 7028 11116 7140 11172
rect 6972 11078 7028 11116
rect 5068 10836 5124 10846
rect 5068 10742 5124 10780
rect 4620 10498 4788 10500
rect 4620 10446 4622 10498
rect 4674 10446 4788 10498
rect 4620 10444 4788 10446
rect 4620 10434 4676 10444
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 7084 10164 7140 11116
rect 7196 10164 7252 10174
rect 7084 10108 7196 10164
rect 7196 10098 7252 10108
rect 4284 9996 4788 10052
rect 4060 9044 4116 9054
rect 4172 9044 4228 9772
rect 4732 9154 4788 9996
rect 6972 9828 7028 9838
rect 6972 9734 7028 9772
rect 4732 9102 4734 9154
rect 4786 9102 4788 9154
rect 4732 9090 4788 9102
rect 7308 9266 7364 12012
rect 7868 12002 7924 12012
rect 7868 11508 7924 11518
rect 7868 11414 7924 11452
rect 7756 10836 7812 10846
rect 7756 9938 7812 10780
rect 7756 9886 7758 9938
rect 7810 9886 7812 9938
rect 7756 9874 7812 9886
rect 7308 9214 7310 9266
rect 7362 9214 7364 9266
rect 4060 9042 4228 9044
rect 4060 8990 4062 9042
rect 4114 8990 4228 9042
rect 4060 8988 4228 8990
rect 4060 8978 4116 8988
rect 6860 8932 6916 8942
rect 7196 8932 7252 8942
rect 6860 8930 7252 8932
rect 6860 8878 6862 8930
rect 6914 8878 7198 8930
rect 7250 8878 7252 8930
rect 6860 8876 7252 8878
rect 6860 8866 6916 8876
rect 7196 8866 7252 8876
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 7308 8148 7364 9214
rect 7644 9828 7700 9838
rect 7644 9268 7700 9772
rect 7756 9268 7812 9278
rect 7644 9212 7756 9268
rect 7308 8082 7364 8092
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 7756 6690 7812 9212
rect 7980 8428 8036 13468
rect 8092 12178 8148 13468
rect 8316 13188 8372 15372
rect 8652 15316 8708 15596
rect 9548 15540 9604 20412
rect 9660 20402 9716 20412
rect 9884 20242 9940 20972
rect 9996 20802 10052 21196
rect 9996 20750 9998 20802
rect 10050 20750 10052 20802
rect 9996 20738 10052 20750
rect 10220 20802 10276 21308
rect 10332 21028 10388 21420
rect 10444 21028 10500 21038
rect 10332 21026 10500 21028
rect 10332 20974 10446 21026
rect 10498 20974 10500 21026
rect 10332 20972 10500 20974
rect 10444 20962 10500 20972
rect 10556 21028 10612 22988
rect 10556 20962 10612 20972
rect 10220 20750 10222 20802
rect 10274 20750 10276 20802
rect 10220 20738 10276 20750
rect 10556 20802 10612 20814
rect 10556 20750 10558 20802
rect 10610 20750 10612 20802
rect 9884 20190 9886 20242
rect 9938 20190 9940 20242
rect 9884 20178 9940 20190
rect 10108 20018 10164 20030
rect 10108 19966 10110 20018
rect 10162 19966 10164 20018
rect 9772 19908 9828 19918
rect 9772 19814 9828 19852
rect 10108 19796 10164 19966
rect 10108 19730 10164 19740
rect 10108 19124 10164 19134
rect 10108 19030 10164 19068
rect 10444 19012 10500 19022
rect 10444 18918 10500 18956
rect 10556 17220 10612 20750
rect 11004 20804 11060 25228
rect 11116 25282 11172 25294
rect 11116 25230 11118 25282
rect 11170 25230 11172 25282
rect 11116 24948 11172 25230
rect 11116 24882 11172 24892
rect 11116 24722 11172 24734
rect 11116 24670 11118 24722
rect 11170 24670 11172 24722
rect 11116 24612 11172 24670
rect 11564 24724 11620 25454
rect 11564 24658 11620 24668
rect 11116 24546 11172 24556
rect 11676 24612 11732 26908
rect 12236 26964 12292 27002
rect 12236 26898 12292 26908
rect 15148 25620 15204 32284
rect 15596 30994 15652 31006
rect 15596 30942 15598 30994
rect 15650 30942 15652 30994
rect 15596 30772 15652 30942
rect 16156 30994 16212 31006
rect 16156 30942 16158 30994
rect 16210 30942 16212 30994
rect 16156 30884 16212 30942
rect 16156 30818 16212 30828
rect 16268 30882 16324 30894
rect 16268 30830 16270 30882
rect 16322 30830 16324 30882
rect 15596 30706 15652 30716
rect 16268 30322 16324 30830
rect 16268 30270 16270 30322
rect 16322 30270 16324 30322
rect 16268 30258 16324 30270
rect 16380 30210 16436 32284
rect 16380 30158 16382 30210
rect 16434 30158 16436 30210
rect 16380 30146 16436 30158
rect 16268 29986 16324 29998
rect 16268 29934 16270 29986
rect 16322 29934 16324 29986
rect 15372 29426 15428 29438
rect 15372 29374 15374 29426
rect 15426 29374 15428 29426
rect 15372 29204 15428 29374
rect 15372 29138 15428 29148
rect 15484 29314 15540 29326
rect 15484 29262 15486 29314
rect 15538 29262 15540 29314
rect 15484 27972 15540 29262
rect 15932 29314 15988 29326
rect 15932 29262 15934 29314
rect 15986 29262 15988 29314
rect 15932 29204 15988 29262
rect 15932 29138 15988 29148
rect 15484 27906 15540 27916
rect 16156 27860 16212 27870
rect 16156 27766 16212 27804
rect 15148 25554 15204 25564
rect 16268 25506 16324 29934
rect 16268 25454 16270 25506
rect 16322 25454 16324 25506
rect 16268 25442 16324 25454
rect 11900 25284 11956 25294
rect 11900 25190 11956 25228
rect 11900 24948 11956 24958
rect 11900 24834 11956 24892
rect 11900 24782 11902 24834
rect 11954 24782 11956 24834
rect 11900 24770 11956 24782
rect 14476 24724 14532 24734
rect 14476 24630 14532 24668
rect 16156 24724 16212 24734
rect 16156 24630 16212 24668
rect 11676 24546 11732 24556
rect 12348 24612 12404 24622
rect 12348 23380 12404 24556
rect 14028 24612 14084 24622
rect 14364 24612 14420 24622
rect 14028 24610 14420 24612
rect 14028 24558 14030 24610
rect 14082 24558 14366 24610
rect 14418 24558 14420 24610
rect 14028 24556 14420 24558
rect 14028 24546 14084 24556
rect 14364 24546 14420 24556
rect 15708 23940 15764 23950
rect 15372 23828 15428 23838
rect 15372 23734 15428 23772
rect 12348 23378 12740 23380
rect 12348 23326 12350 23378
rect 12402 23326 12740 23378
rect 12348 23324 12740 23326
rect 12348 23314 12404 23324
rect 12684 23154 12740 23324
rect 12684 23102 12686 23154
rect 12738 23102 12740 23154
rect 11340 23042 11396 23054
rect 11340 22990 11342 23042
rect 11394 22990 11396 23042
rect 11340 21700 11396 22990
rect 12684 21812 12740 23102
rect 13468 23044 13524 23054
rect 13468 22950 13524 22988
rect 15596 23044 15652 23054
rect 15708 23044 15764 23884
rect 15596 23042 15764 23044
rect 15596 22990 15598 23042
rect 15650 22990 15764 23042
rect 15596 22988 15764 22990
rect 15596 22978 15652 22988
rect 12684 21746 12740 21756
rect 13468 21810 13524 21822
rect 13468 21758 13470 21810
rect 13522 21758 13524 21810
rect 11340 21634 11396 21644
rect 13468 21700 13524 21758
rect 14028 21812 14084 21822
rect 14028 21718 14084 21756
rect 13468 21634 13524 21644
rect 11004 20738 11060 20748
rect 11228 21474 11284 21486
rect 11228 21422 11230 21474
rect 11282 21422 11284 21474
rect 10780 20580 10836 20590
rect 11228 20580 11284 21422
rect 15036 21474 15092 21486
rect 15036 21422 15038 21474
rect 15090 21422 15092 21474
rect 15036 21364 15092 21422
rect 14588 20916 14644 20926
rect 14140 20914 14644 20916
rect 14140 20862 14590 20914
rect 14642 20862 14644 20914
rect 14140 20860 14644 20862
rect 14140 20802 14196 20860
rect 14588 20850 14644 20860
rect 14140 20750 14142 20802
rect 14194 20750 14196 20802
rect 14140 20738 14196 20750
rect 14812 20804 14868 20814
rect 15036 20804 15092 21308
rect 14812 20802 15092 20804
rect 14812 20750 14814 20802
rect 14866 20750 15092 20802
rect 14812 20748 15092 20750
rect 15596 21474 15652 21486
rect 15596 21422 15598 21474
rect 15650 21422 15652 21474
rect 15596 20804 15652 21422
rect 15596 20802 15764 20804
rect 15596 20750 15598 20802
rect 15650 20750 15764 20802
rect 15596 20748 15764 20750
rect 14812 20738 14868 20748
rect 15596 20738 15652 20748
rect 13804 20692 13860 20702
rect 14476 20692 14532 20702
rect 13804 20598 13860 20636
rect 14364 20690 14532 20692
rect 14364 20638 14478 20690
rect 14530 20638 14532 20690
rect 14364 20636 14532 20638
rect 10780 20578 11284 20580
rect 10780 20526 10782 20578
rect 10834 20526 11284 20578
rect 10780 20524 11284 20526
rect 10780 20514 10836 20524
rect 12012 19908 12068 19918
rect 11116 19796 11172 19806
rect 11004 19234 11060 19246
rect 11004 19182 11006 19234
rect 11058 19182 11060 19234
rect 11004 19012 11060 19182
rect 11004 18946 11060 18956
rect 10220 16996 10276 17006
rect 10108 16940 10220 16996
rect 9660 16884 9716 16894
rect 9660 16790 9716 16828
rect 9884 16548 9940 16558
rect 9884 16098 9940 16492
rect 9884 16046 9886 16098
rect 9938 16046 9940 16098
rect 9660 15540 9716 15550
rect 8876 15538 9716 15540
rect 8876 15486 9662 15538
rect 9714 15486 9716 15538
rect 8876 15484 9716 15486
rect 8764 15428 8820 15438
rect 8764 15334 8820 15372
rect 8876 15426 8932 15484
rect 8876 15374 8878 15426
rect 8930 15374 8932 15426
rect 8876 15362 8932 15374
rect 8652 15148 8708 15260
rect 8540 15092 8708 15148
rect 9436 15204 9492 15484
rect 9660 15474 9716 15484
rect 9436 15138 9492 15148
rect 9548 15316 9604 15326
rect 8540 14306 8596 15092
rect 8540 14254 8542 14306
rect 8594 14254 8596 14306
rect 8540 14196 8596 14254
rect 8540 14140 9156 14196
rect 8316 13122 8372 13132
rect 8092 12126 8094 12178
rect 8146 12126 8148 12178
rect 8092 12114 8148 12126
rect 8316 11956 8372 11966
rect 8316 11862 8372 11900
rect 8764 11954 8820 11966
rect 8764 11902 8766 11954
rect 8818 11902 8820 11954
rect 8204 11508 8260 11518
rect 8204 11394 8260 11452
rect 8204 11342 8206 11394
rect 8258 11342 8260 11394
rect 8204 11330 8260 11342
rect 8540 11394 8596 11406
rect 8540 11342 8542 11394
rect 8594 11342 8596 11394
rect 8540 11060 8596 11342
rect 8764 11394 8820 11902
rect 8764 11342 8766 11394
rect 8818 11342 8820 11394
rect 8764 11330 8820 11342
rect 8652 11284 8708 11294
rect 8652 11190 8708 11228
rect 8988 11170 9044 11182
rect 8988 11118 8990 11170
rect 9042 11118 9044 11170
rect 8988 11060 9044 11118
rect 8540 11004 9044 11060
rect 7868 8372 8036 8428
rect 7868 8260 7924 8372
rect 7868 8166 7924 8204
rect 8540 8260 8596 8270
rect 8988 8260 9044 8270
rect 8540 8258 8708 8260
rect 8540 8206 8542 8258
rect 8594 8206 8708 8258
rect 8540 8204 8708 8206
rect 8540 8194 8596 8204
rect 8652 8146 8708 8204
rect 8988 8166 9044 8204
rect 8652 8094 8654 8146
rect 8706 8094 8708 8146
rect 8652 8082 8708 8094
rect 8876 8148 8932 8158
rect 8876 8054 8932 8092
rect 7980 8034 8036 8046
rect 7980 7982 7982 8034
rect 8034 7982 8036 8034
rect 7980 7588 8036 7982
rect 8092 8036 8148 8046
rect 8092 7942 8148 7980
rect 8316 7700 8372 7710
rect 8316 7606 8372 7644
rect 8988 7700 9044 7710
rect 9100 7700 9156 14140
rect 9548 13970 9604 15260
rect 9884 15316 9940 16046
rect 10108 16098 10164 16940
rect 10220 16930 10276 16940
rect 10332 16772 10388 16782
rect 10108 16046 10110 16098
rect 10162 16046 10164 16098
rect 10108 16034 10164 16046
rect 10220 16770 10388 16772
rect 10220 16718 10334 16770
rect 10386 16718 10388 16770
rect 10220 16716 10388 16718
rect 10220 15874 10276 16716
rect 10332 16706 10388 16716
rect 10220 15822 10222 15874
rect 10274 15822 10276 15874
rect 10220 15810 10276 15822
rect 10444 16322 10500 16334
rect 10444 16270 10446 16322
rect 10498 16270 10500 16322
rect 10444 15764 10500 16270
rect 10556 16098 10612 17164
rect 10556 16046 10558 16098
rect 10610 16046 10612 16098
rect 10556 16034 10612 16046
rect 10444 15708 11060 15764
rect 9884 15250 9940 15260
rect 9548 13918 9550 13970
rect 9602 13918 9604 13970
rect 9548 12292 9604 13918
rect 9772 15204 9828 15214
rect 9772 13972 9828 15148
rect 10444 15092 10500 15102
rect 10444 14530 10500 15036
rect 10444 14478 10446 14530
rect 10498 14478 10500 14530
rect 10444 14466 10500 14478
rect 11004 14420 11060 15708
rect 11116 15092 11172 19740
rect 11452 19460 11508 19470
rect 11452 19366 11508 19404
rect 11228 19348 11284 19358
rect 11228 19254 11284 19292
rect 12012 19348 12068 19852
rect 12012 19254 12068 19292
rect 11564 19122 11620 19134
rect 11564 19070 11566 19122
rect 11618 19070 11620 19122
rect 11564 17108 11620 19070
rect 14364 19124 14420 20636
rect 14476 20626 14532 20636
rect 15260 20692 15316 20702
rect 15260 20598 15316 20636
rect 14364 19058 14420 19068
rect 14476 20132 14532 20142
rect 11564 17042 11620 17052
rect 11900 18450 11956 18462
rect 11900 18398 11902 18450
rect 11954 18398 11956 18450
rect 11676 16996 11732 17006
rect 11676 16322 11732 16940
rect 11676 16270 11678 16322
rect 11730 16270 11732 16322
rect 11676 16258 11732 16270
rect 11900 16884 11956 18398
rect 12572 18338 12628 18350
rect 12572 18286 12574 18338
rect 12626 18286 12628 18338
rect 11788 16100 11844 16110
rect 11788 16006 11844 16044
rect 11900 15876 11956 16828
rect 12348 17108 12404 17118
rect 12572 17108 12628 18286
rect 13468 17220 13524 17230
rect 12908 17108 12964 17118
rect 12572 17106 12964 17108
rect 12572 17054 12910 17106
rect 12962 17054 12964 17106
rect 12572 17052 12964 17054
rect 11900 15810 11956 15820
rect 12124 16324 12180 16334
rect 11116 15026 11172 15036
rect 12124 15538 12180 16268
rect 12124 15486 12126 15538
rect 12178 15486 12180 15538
rect 11340 14532 11396 14542
rect 11340 14438 11396 14476
rect 12012 14532 12068 14542
rect 12124 14532 12180 15486
rect 12348 15540 12404 17052
rect 12908 17042 12964 17052
rect 13132 17108 13188 17118
rect 13020 16996 13076 17006
rect 13020 16902 13076 16940
rect 12796 16882 12852 16894
rect 12796 16830 12798 16882
rect 12850 16830 12852 16882
rect 12460 16770 12516 16782
rect 12460 16718 12462 16770
rect 12514 16718 12516 16770
rect 12460 16100 12516 16718
rect 12796 16772 12852 16830
rect 13132 16772 13188 17052
rect 13244 16884 13300 16894
rect 13244 16790 13300 16828
rect 13468 16882 13524 17164
rect 13468 16830 13470 16882
rect 13522 16830 13524 16882
rect 13468 16818 13524 16830
rect 14476 16994 14532 20076
rect 15148 20130 15204 20142
rect 15148 20078 15150 20130
rect 15202 20078 15204 20130
rect 14924 20020 14980 20030
rect 14924 19926 14980 19964
rect 15148 19796 15204 20078
rect 15484 20020 15540 20030
rect 15484 19926 15540 19964
rect 15148 19730 15204 19740
rect 15372 19348 15428 19358
rect 15708 19348 15764 20748
rect 16380 20692 16436 20702
rect 16380 20598 16436 20636
rect 15820 20132 15876 20142
rect 15820 20038 15876 20076
rect 16492 20132 16548 32396
rect 16604 31892 16660 32508
rect 16828 32452 16884 32462
rect 16940 32452 16996 32462
rect 16828 32450 16940 32452
rect 16828 32398 16830 32450
rect 16882 32398 16940 32450
rect 16828 32396 16940 32398
rect 16828 32386 16884 32396
rect 16604 31826 16660 31836
rect 16716 30884 16772 30894
rect 16716 30790 16772 30828
rect 16828 29316 16884 29326
rect 16828 28642 16884 29260
rect 16828 28590 16830 28642
rect 16882 28590 16884 28642
rect 16828 28578 16884 28590
rect 16604 28084 16660 28094
rect 16604 25394 16660 28028
rect 16716 27860 16772 27870
rect 16716 27766 16772 27804
rect 16828 27748 16884 27758
rect 16828 27654 16884 27692
rect 16604 25342 16606 25394
rect 16658 25342 16660 25394
rect 16604 25330 16660 25342
rect 16828 25396 16884 25406
rect 16716 24948 16772 24958
rect 16716 24722 16772 24892
rect 16828 24834 16884 25340
rect 16828 24782 16830 24834
rect 16882 24782 16884 24834
rect 16828 24770 16884 24782
rect 16716 24670 16718 24722
rect 16770 24670 16772 24722
rect 16716 24658 16772 24670
rect 16940 21700 16996 32396
rect 17388 29428 17444 38670
rect 17612 38836 17668 38846
rect 17612 38722 17668 38780
rect 17612 38670 17614 38722
rect 17666 38670 17668 38722
rect 17612 38668 17668 38670
rect 17500 38612 17668 38668
rect 17500 30436 17556 38612
rect 17724 37940 17780 39454
rect 18172 38948 18228 38958
rect 17948 38834 18004 38846
rect 17948 38782 17950 38834
rect 18002 38782 18004 38834
rect 17948 38610 18004 38782
rect 17948 38558 17950 38610
rect 18002 38558 18004 38610
rect 17948 38546 18004 38558
rect 17948 38276 18004 38286
rect 18172 38276 18228 38892
rect 17948 38274 18228 38276
rect 17948 38222 17950 38274
rect 18002 38222 18228 38274
rect 17948 38220 18228 38222
rect 19068 38388 19124 38398
rect 17948 38210 18004 38220
rect 18060 38052 18116 38062
rect 18060 37958 18116 37996
rect 18284 38050 18340 38062
rect 18508 38052 18564 38062
rect 18284 37998 18286 38050
rect 18338 37998 18340 38050
rect 17724 37874 17780 37884
rect 18284 36596 18340 37998
rect 18284 36530 18340 36540
rect 18396 38050 18564 38052
rect 18396 37998 18510 38050
rect 18562 37998 18564 38050
rect 18396 37996 18564 37998
rect 18396 36594 18452 37996
rect 18508 37986 18564 37996
rect 18620 38050 18676 38062
rect 18620 37998 18622 38050
rect 18674 37998 18676 38050
rect 18508 37380 18564 37390
rect 18620 37380 18676 37998
rect 19068 37938 19124 38332
rect 19068 37886 19070 37938
rect 19122 37886 19124 37938
rect 19068 37874 19124 37886
rect 18508 37378 18676 37380
rect 18508 37326 18510 37378
rect 18562 37326 18676 37378
rect 18508 37324 18676 37326
rect 18508 37314 18564 37324
rect 19068 37268 19124 37278
rect 19068 37174 19124 37212
rect 18396 36542 18398 36594
rect 18450 36542 18452 36594
rect 18396 36530 18452 36542
rect 18732 36596 18788 36606
rect 18732 36502 18788 36540
rect 17724 36484 17780 36494
rect 17724 36390 17780 36428
rect 18172 36482 18228 36494
rect 18172 36430 18174 36482
rect 18226 36430 18228 36482
rect 17948 34020 18004 34030
rect 17948 33346 18004 33964
rect 17948 33294 17950 33346
rect 18002 33294 18004 33346
rect 17836 32562 17892 32574
rect 17836 32510 17838 32562
rect 17890 32510 17892 32562
rect 17724 32452 17780 32462
rect 17836 32452 17892 32510
rect 17780 32396 17892 32452
rect 17724 32386 17780 32396
rect 17836 31780 17892 31790
rect 17948 31780 18004 33294
rect 17836 31778 18004 31780
rect 17836 31726 17838 31778
rect 17890 31726 18004 31778
rect 17836 31724 18004 31726
rect 17836 31556 17892 31724
rect 17836 31490 17892 31500
rect 17948 30996 18004 31006
rect 17948 30902 18004 30940
rect 18172 30882 18228 36430
rect 18844 36482 18900 36494
rect 18844 36430 18846 36482
rect 18898 36430 18900 36482
rect 18508 35252 18564 35262
rect 18508 34914 18564 35196
rect 18508 34862 18510 34914
rect 18562 34862 18564 34914
rect 18508 34850 18564 34862
rect 18844 34914 18900 36430
rect 19180 36484 19236 36494
rect 19180 36390 19236 36428
rect 19292 35588 19348 39566
rect 19404 39506 19460 39518
rect 19404 39454 19406 39506
rect 19458 39454 19460 39506
rect 19404 38668 19460 39454
rect 19516 39058 19572 41580
rect 19628 40962 19684 40974
rect 19628 40910 19630 40962
rect 19682 40910 19684 40962
rect 19628 40404 19684 40910
rect 19836 40796 20100 40806
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 19836 40730 20100 40740
rect 19740 40516 19796 40526
rect 19740 40422 19796 40460
rect 19628 40338 19684 40348
rect 19836 39228 20100 39238
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 19836 39162 20100 39172
rect 19516 39006 19518 39058
rect 19570 39006 19572 39058
rect 19516 38994 19572 39006
rect 19740 38948 19796 38958
rect 19740 38854 19796 38892
rect 19852 38834 19908 38846
rect 19852 38782 19854 38834
rect 19906 38782 19908 38834
rect 19852 38668 19908 38782
rect 20188 38722 20244 38734
rect 20188 38670 20190 38722
rect 20242 38670 20244 38722
rect 19404 38612 19684 38668
rect 19852 38612 20020 38668
rect 19628 38050 19684 38612
rect 19964 38162 20020 38612
rect 19964 38110 19966 38162
rect 20018 38110 20020 38162
rect 19964 38098 20020 38110
rect 19628 37998 19630 38050
rect 19682 37998 19684 38050
rect 19628 37986 19684 37998
rect 20188 38050 20244 38670
rect 20188 37998 20190 38050
rect 20242 37998 20244 38050
rect 20188 37986 20244 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 19404 37156 19460 37166
rect 20076 37156 20132 37166
rect 19404 37154 20132 37156
rect 19404 37102 19406 37154
rect 19458 37102 20078 37154
rect 20130 37102 20132 37154
rect 19404 37100 20132 37102
rect 19404 37090 19460 37100
rect 20076 36372 20132 37100
rect 20076 36306 20132 36316
rect 20188 36258 20244 36270
rect 20188 36206 20190 36258
rect 20242 36206 20244 36258
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19292 35522 19348 35532
rect 18844 34862 18846 34914
rect 18898 34862 18900 34914
rect 18844 34692 18900 34862
rect 18844 34626 18900 34636
rect 18956 34802 19012 34814
rect 18956 34750 18958 34802
rect 19010 34750 19012 34802
rect 18732 34244 18788 34254
rect 18396 34188 18732 34244
rect 18284 34018 18340 34030
rect 18284 33966 18286 34018
rect 18338 33966 18340 34018
rect 18284 32900 18340 33966
rect 18284 32834 18340 32844
rect 18396 32562 18452 34188
rect 18732 34150 18788 34188
rect 18956 33572 19012 34750
rect 19404 34692 19460 34702
rect 19404 34598 19460 34636
rect 20188 34692 20244 36206
rect 20188 34626 20244 34636
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19180 34020 19236 34030
rect 19180 33926 19236 33964
rect 18956 33506 19012 33516
rect 19628 33460 19684 33470
rect 18844 33346 18900 33358
rect 18844 33294 18846 33346
rect 18898 33294 18900 33346
rect 18844 32900 18900 33294
rect 19404 33348 19460 33358
rect 19404 33254 19460 33292
rect 18844 32834 18900 32844
rect 19516 33234 19572 33246
rect 19516 33182 19518 33234
rect 19570 33182 19572 33234
rect 19068 32786 19124 32798
rect 19068 32734 19070 32786
rect 19122 32734 19124 32786
rect 18956 32674 19012 32686
rect 18956 32622 18958 32674
rect 19010 32622 19012 32674
rect 18396 32510 18398 32562
rect 18450 32510 18452 32562
rect 18396 32498 18452 32510
rect 18508 32564 18564 32574
rect 18844 32564 18900 32574
rect 18508 32562 18900 32564
rect 18508 32510 18510 32562
rect 18562 32510 18846 32562
rect 18898 32510 18900 32562
rect 18508 32508 18900 32510
rect 18508 32498 18564 32508
rect 18844 32498 18900 32508
rect 18172 30830 18174 30882
rect 18226 30830 18228 30882
rect 17500 30380 17668 30436
rect 17500 29428 17556 29438
rect 17388 29372 17500 29428
rect 17500 29334 17556 29372
rect 17276 28644 17332 28654
rect 17276 28550 17332 28588
rect 17388 28530 17444 28542
rect 17388 28478 17390 28530
rect 17442 28478 17444 28530
rect 17164 27860 17220 27870
rect 17164 27636 17220 27804
rect 17388 27858 17444 28478
rect 17500 27972 17556 27982
rect 17500 27878 17556 27916
rect 17388 27806 17390 27858
rect 17442 27806 17444 27858
rect 17388 27794 17444 27806
rect 17164 27186 17220 27580
rect 17164 27134 17166 27186
rect 17218 27134 17220 27186
rect 17164 27122 17220 27134
rect 17612 26908 17668 30380
rect 17724 30212 17780 30222
rect 17724 29426 17780 30156
rect 18172 30100 18228 30830
rect 18172 30034 18228 30044
rect 18508 31892 18564 31902
rect 18508 30996 18564 31836
rect 18620 31108 18676 31118
rect 18956 31108 19012 32622
rect 19068 32676 19124 32734
rect 19068 32610 19124 32620
rect 19516 32564 19572 33182
rect 19516 32498 19572 32508
rect 18620 31106 19012 31108
rect 18620 31054 18622 31106
rect 18674 31054 19012 31106
rect 18620 31052 19012 31054
rect 19628 31890 19684 33404
rect 19964 33348 20020 33358
rect 19964 33254 20020 33292
rect 20300 33012 20356 43652
rect 20748 43652 20804 43662
rect 21084 43652 21140 43662
rect 20804 43650 21140 43652
rect 20804 43598 21086 43650
rect 21138 43598 21140 43650
rect 20804 43596 21140 43598
rect 20748 43558 20804 43596
rect 21084 43586 21140 43596
rect 20412 43540 20468 43550
rect 20412 43446 20468 43484
rect 22652 41746 22708 44492
rect 22764 43876 22820 50316
rect 23996 50036 24052 50430
rect 24108 50484 24164 50494
rect 24108 50390 24164 50428
rect 24556 50484 24612 50494
rect 25004 50482 25060 50494
rect 25004 50430 25006 50482
rect 25058 50430 25060 50482
rect 25004 50428 25060 50430
rect 24556 50390 24612 50428
rect 24892 50372 25060 50428
rect 25116 50484 25172 50494
rect 25900 50484 25956 50494
rect 25116 50390 25172 50428
rect 25788 50372 25956 50428
rect 24108 50036 24164 50046
rect 23996 50034 24164 50036
rect 23996 49982 24110 50034
rect 24162 49982 24164 50034
rect 23996 49980 24164 49982
rect 24108 49970 24164 49980
rect 24556 49812 24612 49822
rect 22876 49700 22932 49710
rect 23212 49700 23268 49710
rect 22876 49698 23212 49700
rect 22876 49646 22878 49698
rect 22930 49646 23212 49698
rect 22876 49644 23212 49646
rect 22876 49634 22932 49644
rect 23212 49606 23268 49644
rect 23436 49586 23492 49598
rect 23436 49534 23438 49586
rect 23490 49534 23492 49586
rect 23436 48580 23492 49534
rect 23436 48514 23492 48524
rect 23660 49586 23716 49598
rect 23660 49534 23662 49586
rect 23714 49534 23716 49586
rect 23100 48244 23156 48254
rect 23100 48150 23156 48188
rect 23660 48132 23716 49534
rect 24444 48692 24500 48702
rect 24332 48356 24388 48366
rect 23996 48242 24052 48254
rect 23996 48190 23998 48242
rect 24050 48190 24052 48242
rect 23996 48132 24052 48190
rect 23660 48076 24052 48132
rect 23772 47346 23828 48076
rect 24220 48018 24276 48030
rect 24220 47966 24222 48018
rect 24274 47966 24276 48018
rect 24108 47572 24164 47582
rect 24108 47478 24164 47516
rect 23772 47294 23774 47346
rect 23826 47294 23828 47346
rect 23436 46788 23492 46798
rect 23436 45892 23492 46732
rect 23436 45826 23492 45836
rect 22876 45444 22932 45454
rect 22876 45330 22932 45388
rect 23772 45444 23828 47294
rect 23996 47236 24052 47246
rect 24220 47236 24276 47966
rect 23996 47234 24276 47236
rect 23996 47182 23998 47234
rect 24050 47182 24276 47234
rect 23996 47180 24276 47182
rect 23996 46788 24052 47180
rect 23996 46722 24052 46732
rect 24332 45778 24388 48300
rect 24444 48242 24500 48636
rect 24556 48354 24612 49756
rect 24556 48302 24558 48354
rect 24610 48302 24612 48354
rect 24556 48290 24612 48302
rect 24892 49700 24948 50372
rect 24444 48190 24446 48242
rect 24498 48190 24500 48242
rect 24444 48178 24500 48190
rect 24444 47346 24500 47358
rect 24444 47294 24446 47346
rect 24498 47294 24500 47346
rect 24444 46788 24500 47294
rect 24780 47348 24836 47358
rect 24892 47348 24948 49644
rect 25228 49810 25284 49822
rect 25228 49758 25230 49810
rect 25282 49758 25284 49810
rect 25228 49028 25284 49758
rect 25452 49812 25508 49822
rect 25452 49718 25508 49756
rect 25676 49810 25732 49822
rect 25676 49758 25678 49810
rect 25730 49758 25732 49810
rect 25564 49700 25620 49710
rect 25564 49606 25620 49644
rect 25284 48972 25396 49028
rect 25228 48962 25284 48972
rect 24780 47346 24948 47348
rect 24780 47294 24782 47346
rect 24834 47294 24948 47346
rect 24780 47292 24948 47294
rect 24780 47282 24836 47292
rect 24444 46722 24500 46732
rect 24668 46676 24724 46686
rect 24668 46674 24836 46676
rect 24668 46622 24670 46674
rect 24722 46622 24836 46674
rect 24668 46620 24836 46622
rect 24668 46610 24724 46620
rect 24332 45726 24334 45778
rect 24386 45726 24388 45778
rect 24332 45714 24388 45726
rect 23772 45378 23828 45388
rect 23996 45666 24052 45678
rect 23996 45614 23998 45666
rect 24050 45614 24052 45666
rect 22876 45278 22878 45330
rect 22930 45278 22932 45330
rect 22876 45266 22932 45278
rect 23212 45332 23268 45342
rect 23212 45238 23268 45276
rect 23436 45106 23492 45118
rect 23436 45054 23438 45106
rect 23490 45054 23492 45106
rect 23436 44884 23492 45054
rect 23996 44996 24052 45614
rect 24668 45668 24724 45678
rect 23996 44930 24052 44940
rect 24556 44996 24612 45006
rect 24668 44996 24724 45612
rect 24612 44940 24724 44996
rect 24556 44902 24612 44940
rect 22876 44324 22932 44334
rect 23436 44324 23492 44828
rect 24668 44772 24724 44940
rect 24668 44706 24724 44716
rect 24780 45556 24836 46620
rect 22876 44322 23492 44324
rect 22876 44270 22878 44322
rect 22930 44270 23438 44322
rect 23490 44270 23492 44322
rect 22876 44268 23492 44270
rect 22876 44258 22932 44268
rect 23436 44258 23492 44268
rect 23212 44100 23268 44110
rect 23436 44100 23492 44110
rect 23212 44006 23268 44044
rect 23324 44044 23436 44100
rect 22764 43820 22932 43876
rect 22652 41694 22654 41746
rect 22706 41694 22708 41746
rect 22652 41682 22708 41694
rect 22204 41188 22260 41198
rect 22764 41188 22820 41198
rect 21868 41186 22820 41188
rect 21868 41134 22206 41186
rect 22258 41134 22766 41186
rect 22818 41134 22820 41186
rect 21868 41132 22820 41134
rect 20860 40292 20916 40302
rect 20860 38834 20916 40236
rect 21868 40292 21924 41132
rect 22204 41122 22260 41132
rect 22764 41122 22820 41132
rect 22428 40964 22484 40974
rect 22428 40870 22484 40908
rect 21868 40198 21924 40236
rect 22092 40740 22148 40750
rect 20860 38782 20862 38834
rect 20914 38782 20916 38834
rect 20860 38770 20916 38782
rect 21644 38834 21700 38846
rect 21644 38782 21646 38834
rect 21698 38782 21700 38834
rect 21084 38722 21140 38734
rect 21084 38670 21086 38722
rect 21138 38670 21140 38722
rect 21084 38668 21140 38670
rect 21084 38612 21476 38668
rect 20636 37940 20692 37950
rect 20636 37846 20692 37884
rect 21420 37828 21476 38612
rect 21420 37826 21588 37828
rect 21420 37774 21422 37826
rect 21474 37774 21588 37826
rect 21420 37772 21588 37774
rect 21420 37762 21476 37772
rect 20636 36484 20692 36494
rect 20524 36428 20636 36484
rect 20524 34130 20580 36428
rect 20636 36418 20692 36428
rect 20748 35588 20804 35598
rect 20524 34078 20526 34130
rect 20578 34078 20580 34130
rect 20524 33684 20580 34078
rect 20524 33618 20580 33628
rect 20636 34916 20692 34926
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20300 32946 20356 32956
rect 20412 33572 20468 33582
rect 19836 32890 20100 32900
rect 20412 32674 20468 33516
rect 20636 33348 20692 34860
rect 20412 32622 20414 32674
rect 20466 32622 20468 32674
rect 20412 32610 20468 32622
rect 20524 33292 20692 33348
rect 20748 34020 20804 35532
rect 20524 33234 20580 33292
rect 20524 33182 20526 33234
rect 20578 33182 20580 33234
rect 19852 32564 19908 32574
rect 19852 32470 19908 32508
rect 19628 31838 19630 31890
rect 19682 31838 19684 31890
rect 18620 31042 18676 31052
rect 17724 29374 17726 29426
rect 17778 29374 17780 29426
rect 17724 29362 17780 29374
rect 17836 29316 17892 29326
rect 17836 28644 17892 29260
rect 17836 28550 17892 28588
rect 18396 29314 18452 29326
rect 18396 29262 18398 29314
rect 18450 29262 18452 29314
rect 18396 27972 18452 29262
rect 18396 27906 18452 27916
rect 17500 26852 17668 26908
rect 16940 21634 16996 21644
rect 17052 25618 17108 25630
rect 17052 25566 17054 25618
rect 17106 25566 17108 25618
rect 16492 20066 16548 20076
rect 16716 20692 16772 20702
rect 16156 20020 16212 20030
rect 16156 19908 16212 19964
rect 16604 19908 16660 19918
rect 16156 19906 16660 19908
rect 16156 19854 16606 19906
rect 16658 19854 16660 19906
rect 16156 19852 16660 19854
rect 16604 19796 16660 19852
rect 16604 19730 16660 19740
rect 15148 19346 15764 19348
rect 15148 19294 15374 19346
rect 15426 19294 15764 19346
rect 15148 19292 15764 19294
rect 15148 18674 15204 19292
rect 15372 19282 15428 19292
rect 15708 19234 15764 19292
rect 15708 19182 15710 19234
rect 15762 19182 15764 19234
rect 15708 19170 15764 19182
rect 16492 19124 16548 19134
rect 16492 19122 16660 19124
rect 16492 19070 16494 19122
rect 16546 19070 16660 19122
rect 16492 19068 16660 19070
rect 16492 19058 16548 19068
rect 15148 18622 15150 18674
rect 15202 18622 15204 18674
rect 14700 18338 14756 18350
rect 14700 18286 14702 18338
rect 14754 18286 14756 18338
rect 14700 17556 14756 18286
rect 14700 17490 14756 17500
rect 14812 17780 14868 17790
rect 15148 17780 15204 18622
rect 14476 16942 14478 16994
rect 14530 16942 14532 16994
rect 12796 16716 13188 16772
rect 12460 16034 12516 16044
rect 12684 15876 12740 15886
rect 12684 15782 12740 15820
rect 12796 15540 12852 15550
rect 12348 15538 12852 15540
rect 12348 15486 12798 15538
rect 12850 15486 12852 15538
rect 12348 15484 12852 15486
rect 12348 15314 12404 15484
rect 12796 15474 12852 15484
rect 12348 15262 12350 15314
rect 12402 15262 12404 15314
rect 12348 15250 12404 15262
rect 12908 15148 12964 16716
rect 13132 15428 13188 15438
rect 13132 15334 13188 15372
rect 14364 15428 14420 15438
rect 12068 14476 12180 14532
rect 12572 15092 12964 15148
rect 14028 15314 14084 15326
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 15204 14084 15262
rect 14028 15138 14084 15148
rect 12012 14438 12068 14476
rect 10892 14418 11060 14420
rect 10892 14366 11006 14418
rect 11058 14366 11060 14418
rect 10892 14364 11060 14366
rect 10220 14308 10276 14318
rect 10220 14214 10276 14252
rect 10332 13972 10388 13982
rect 9772 13970 10724 13972
rect 9772 13918 10334 13970
rect 10386 13918 10724 13970
rect 9772 13916 10724 13918
rect 9772 13746 9828 13916
rect 10332 13906 10388 13916
rect 9772 13694 9774 13746
rect 9826 13694 9828 13746
rect 9772 13682 9828 13694
rect 10668 13524 10724 13916
rect 10668 13186 10724 13468
rect 10668 13134 10670 13186
rect 10722 13134 10724 13186
rect 10668 13122 10724 13134
rect 10780 12738 10836 12750
rect 10780 12686 10782 12738
rect 10834 12686 10836 12738
rect 10668 12404 10724 12414
rect 10556 12402 10724 12404
rect 10556 12350 10670 12402
rect 10722 12350 10724 12402
rect 10556 12348 10724 12350
rect 9884 12292 9940 12302
rect 9604 12290 9940 12292
rect 9604 12238 9886 12290
rect 9938 12238 9940 12290
rect 9604 12236 9940 12238
rect 9548 12226 9604 12236
rect 9884 12226 9940 12236
rect 9212 12180 9268 12190
rect 10108 12180 10164 12190
rect 9212 11282 9268 12124
rect 9996 12124 10108 12180
rect 9212 11230 9214 11282
rect 9266 11230 9268 11282
rect 9212 11218 9268 11230
rect 9324 11284 9380 11294
rect 9324 11190 9380 11228
rect 9884 9940 9940 9950
rect 9996 9940 10052 12124
rect 10108 12086 10164 12124
rect 10332 11956 10388 11966
rect 10332 11862 10388 11900
rect 10556 11284 10612 12348
rect 10668 12338 10724 12348
rect 10668 12180 10724 12190
rect 10780 12180 10836 12686
rect 10668 12178 10836 12180
rect 10668 12126 10670 12178
rect 10722 12126 10836 12178
rect 10668 12124 10836 12126
rect 10668 12114 10724 12124
rect 10892 11284 10948 14364
rect 11004 14354 11060 14364
rect 11676 14306 11732 14318
rect 11676 14254 11678 14306
rect 11730 14254 11732 14306
rect 11676 13748 11732 14254
rect 11676 13682 11732 13692
rect 12124 14308 12180 14318
rect 11564 13524 11620 13534
rect 11004 13076 11060 13086
rect 11004 12962 11060 13020
rect 11564 13074 11620 13468
rect 11564 13022 11566 13074
rect 11618 13022 11620 13074
rect 11564 13010 11620 13022
rect 11900 13076 11956 13086
rect 11900 12982 11956 13020
rect 11004 12910 11006 12962
rect 11058 12910 11060 12962
rect 11004 12898 11060 12910
rect 12124 12964 12180 14252
rect 12572 13970 12628 15092
rect 12572 13918 12574 13970
rect 12626 13918 12628 13970
rect 12572 13906 12628 13918
rect 12124 12290 12180 12908
rect 12124 12238 12126 12290
rect 12178 12238 12180 12290
rect 12124 12226 12180 12238
rect 12348 13748 12404 13758
rect 12236 12066 12292 12078
rect 12236 12014 12238 12066
rect 12290 12014 12292 12066
rect 11004 11284 11060 11294
rect 10556 11228 10836 11284
rect 9884 9938 10052 9940
rect 9884 9886 9886 9938
rect 9938 9886 10052 9938
rect 9884 9884 10052 9886
rect 10668 10724 10724 10734
rect 9884 9874 9940 9884
rect 10332 9602 10388 9614
rect 10332 9550 10334 9602
rect 10386 9550 10388 9602
rect 9884 9268 9940 9278
rect 10332 9268 10388 9550
rect 9940 9212 10388 9268
rect 9884 9042 9940 9212
rect 10668 9154 10724 10668
rect 10780 10388 10836 11228
rect 10948 11282 11060 11284
rect 10948 11230 11006 11282
rect 11058 11230 11060 11282
rect 10948 11228 11060 11230
rect 10892 11190 10948 11228
rect 11004 11218 11060 11228
rect 11676 11284 11732 11294
rect 11340 11172 11396 11182
rect 11676 11172 11732 11228
rect 11340 11170 11732 11172
rect 11340 11118 11342 11170
rect 11394 11118 11732 11170
rect 11340 11116 11732 11118
rect 11340 11106 11396 11116
rect 11004 10948 11060 10958
rect 10892 10836 10948 10846
rect 10892 10742 10948 10780
rect 11004 10610 11060 10892
rect 11676 10722 11732 11116
rect 12124 10948 12180 10958
rect 12012 10836 12068 10846
rect 12012 10742 12068 10780
rect 11676 10670 11678 10722
rect 11730 10670 11732 10722
rect 11676 10658 11732 10670
rect 11004 10558 11006 10610
rect 11058 10558 11060 10610
rect 11004 10546 11060 10558
rect 11452 10610 11508 10622
rect 11452 10558 11454 10610
rect 11506 10558 11508 10610
rect 11452 10500 11508 10558
rect 11452 10434 11508 10444
rect 12124 10610 12180 10892
rect 12124 10558 12126 10610
rect 12178 10558 12180 10610
rect 11116 10388 11172 10398
rect 10780 10386 11172 10388
rect 10780 10334 11118 10386
rect 11170 10334 11172 10386
rect 10780 10332 11172 10334
rect 11116 10322 11172 10332
rect 12012 9940 12068 9950
rect 12124 9940 12180 10558
rect 12236 10386 12292 12014
rect 12348 11956 12404 13692
rect 14364 13748 14420 15372
rect 14364 13186 14420 13692
rect 14476 13412 14532 16942
rect 14588 16884 14644 16894
rect 14588 16790 14644 16828
rect 14812 16882 14868 17724
rect 15036 17724 15204 17780
rect 15708 17780 15764 17790
rect 15036 17332 15092 17724
rect 15708 17686 15764 17724
rect 15148 17556 15204 17566
rect 15148 17462 15204 17500
rect 15260 17444 15316 17454
rect 15260 17442 15652 17444
rect 15260 17390 15262 17442
rect 15314 17390 15652 17442
rect 15260 17388 15652 17390
rect 15260 17378 15316 17388
rect 15036 17276 15204 17332
rect 14812 16830 14814 16882
rect 14866 16830 14868 16882
rect 14812 16818 14868 16830
rect 15036 16658 15092 16670
rect 15036 16606 15038 16658
rect 15090 16606 15092 16658
rect 15036 16324 15092 16606
rect 15036 16258 15092 16268
rect 15148 15876 15204 17276
rect 15260 16882 15316 16894
rect 15260 16830 15262 16882
rect 15314 16830 15316 16882
rect 15260 16322 15316 16830
rect 15260 16270 15262 16322
rect 15314 16270 15316 16322
rect 15260 16258 15316 16270
rect 15372 15988 15428 15998
rect 15484 15988 15540 17388
rect 15596 17108 15652 17388
rect 15596 17052 16100 17108
rect 16044 16994 16100 17052
rect 16604 17106 16660 19068
rect 16604 17054 16606 17106
rect 16658 17054 16660 17106
rect 16604 17042 16660 17054
rect 16044 16942 16046 16994
rect 16098 16942 16100 16994
rect 16044 16930 16100 16942
rect 16716 16996 16772 20636
rect 17052 19460 17108 25566
rect 17500 24948 17556 26852
rect 17724 25620 17780 25630
rect 17612 25396 17668 25406
rect 17612 25302 17668 25340
rect 17500 24854 17556 24892
rect 17724 25284 17780 25564
rect 17724 24050 17780 25228
rect 17724 23998 17726 24050
rect 17778 23998 17780 24050
rect 17724 23986 17780 23998
rect 18060 24722 18116 24734
rect 18060 24670 18062 24722
rect 18114 24670 18116 24722
rect 18060 23940 18116 24670
rect 18396 24610 18452 24622
rect 18396 24558 18398 24610
rect 18450 24558 18452 24610
rect 18396 24388 18452 24558
rect 18396 24322 18452 24332
rect 18060 23874 18116 23884
rect 18508 21476 18564 30940
rect 18844 29428 18900 29438
rect 19628 29428 19684 31838
rect 20300 31556 20356 31566
rect 20300 31462 20356 31500
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 20300 30212 20356 30222
rect 20188 30156 20300 30212
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 18900 29372 19236 29428
rect 18844 29334 18900 29372
rect 19180 28756 19236 29372
rect 19180 28662 19236 28700
rect 19292 29426 19684 29428
rect 19292 29374 19630 29426
rect 19682 29374 19684 29426
rect 19292 29372 19684 29374
rect 19292 28308 19348 29372
rect 19628 29362 19684 29372
rect 19628 28868 19684 28878
rect 19628 28774 19684 28812
rect 19740 28756 19796 28766
rect 19740 28644 19796 28700
rect 19628 28588 19796 28644
rect 19180 28252 19348 28308
rect 19516 28530 19572 28542
rect 19516 28478 19518 28530
rect 19570 28478 19572 28530
rect 18844 28084 18900 28094
rect 18844 27990 18900 28028
rect 19068 27076 19124 27086
rect 19068 26982 19124 27020
rect 18956 26962 19012 26974
rect 18956 26910 18958 26962
rect 19010 26910 19012 26962
rect 18956 26068 19012 26910
rect 19068 26292 19124 26302
rect 19180 26292 19236 28252
rect 19404 27858 19460 27870
rect 19404 27806 19406 27858
rect 19458 27806 19460 27858
rect 19404 27748 19460 27806
rect 19404 27682 19460 27692
rect 19516 27524 19572 28478
rect 19628 28530 19684 28588
rect 19628 28478 19630 28530
rect 19682 28478 19684 28530
rect 19628 28466 19684 28478
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19964 27972 20020 27982
rect 19964 27878 20020 27916
rect 19628 27748 19684 27758
rect 19684 27692 19796 27748
rect 19628 27682 19684 27692
rect 19516 27458 19572 27468
rect 19068 26290 19236 26292
rect 19068 26238 19070 26290
rect 19122 26238 19236 26290
rect 19068 26236 19236 26238
rect 19292 27412 19348 27422
rect 19292 26962 19348 27356
rect 19628 27076 19684 27086
rect 19740 27076 19796 27692
rect 19628 27074 19796 27076
rect 19628 27022 19630 27074
rect 19682 27022 19796 27074
rect 19628 27020 19796 27022
rect 19964 27076 20020 27086
rect 19628 27010 19684 27020
rect 19964 26982 20020 27020
rect 20188 27074 20244 30156
rect 20300 30146 20356 30156
rect 20524 30210 20580 33182
rect 20636 33124 20692 33134
rect 20748 33124 20804 33964
rect 21196 34020 21252 34030
rect 21196 34018 21476 34020
rect 21196 33966 21198 34018
rect 21250 33966 21476 34018
rect 21196 33964 21476 33966
rect 21196 33954 21252 33964
rect 21420 33458 21476 33964
rect 21420 33406 21422 33458
rect 21474 33406 21476 33458
rect 21420 33394 21476 33406
rect 20860 33348 20916 33358
rect 21196 33348 21252 33358
rect 20860 33346 21252 33348
rect 20860 33294 20862 33346
rect 20914 33294 21198 33346
rect 21250 33294 21252 33346
rect 20860 33292 21252 33294
rect 20860 33282 20916 33292
rect 21196 33282 21252 33292
rect 21532 33348 21588 37772
rect 21644 36484 21700 38782
rect 21644 36390 21700 36428
rect 21868 36372 21924 36382
rect 21868 35922 21924 36316
rect 21868 35870 21870 35922
rect 21922 35870 21924 35922
rect 21868 35858 21924 35870
rect 21532 33282 21588 33292
rect 21644 33236 21700 33246
rect 21644 33142 21700 33180
rect 21868 33234 21924 33246
rect 21868 33182 21870 33234
rect 21922 33182 21924 33234
rect 20636 33122 20804 33124
rect 20636 33070 20638 33122
rect 20690 33070 20804 33122
rect 20636 33068 20804 33070
rect 20860 33124 20916 33134
rect 20636 33058 20692 33068
rect 20860 32786 20916 33068
rect 20860 32734 20862 32786
rect 20914 32734 20916 32786
rect 20860 32722 20916 32734
rect 21196 32562 21252 32574
rect 21196 32510 21198 32562
rect 21250 32510 21252 32562
rect 21196 32452 21252 32510
rect 21644 32452 21700 32462
rect 21196 32450 21700 32452
rect 21196 32398 21646 32450
rect 21698 32398 21700 32450
rect 21196 32396 21700 32398
rect 21644 32340 21700 32396
rect 20524 30158 20526 30210
rect 20578 30158 20580 30210
rect 20412 29988 20468 29998
rect 20188 27022 20190 27074
rect 20242 27022 20244 27074
rect 19292 26910 19294 26962
rect 19346 26910 19348 26962
rect 19068 26226 19124 26236
rect 19292 26068 19348 26910
rect 19404 26964 19460 26974
rect 19404 26870 19460 26908
rect 19852 26852 19908 26862
rect 19628 26850 19908 26852
rect 19628 26798 19854 26850
rect 19906 26798 19908 26850
rect 19628 26796 19908 26798
rect 19628 26404 19684 26796
rect 19852 26786 19908 26796
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19740 26404 19796 26414
rect 19628 26402 19796 26404
rect 19628 26350 19742 26402
rect 19794 26350 19796 26402
rect 19628 26348 19796 26350
rect 19740 26338 19796 26348
rect 18956 26012 19348 26068
rect 19180 25506 19236 25518
rect 19180 25454 19182 25506
rect 19234 25454 19236 25506
rect 18956 24836 19012 24846
rect 19180 24836 19236 25454
rect 19292 25172 19348 26012
rect 19852 25508 19908 25518
rect 19852 25414 19908 25452
rect 19516 25282 19572 25294
rect 19516 25230 19518 25282
rect 19570 25230 19572 25282
rect 19292 25116 19460 25172
rect 18956 24834 19236 24836
rect 18956 24782 18958 24834
rect 19010 24782 19236 24834
rect 18956 24780 19236 24782
rect 18956 24770 19012 24780
rect 19292 24388 19348 24398
rect 19292 23378 19348 24332
rect 19292 23326 19294 23378
rect 19346 23326 19348 23378
rect 19292 23314 19348 23326
rect 19180 21476 19236 21486
rect 18508 21474 19236 21476
rect 18508 21422 19182 21474
rect 19234 21422 19236 21474
rect 18508 21420 19236 21422
rect 18508 20916 18564 20926
rect 18508 20822 18564 20860
rect 19068 20802 19124 20814
rect 19068 20750 19070 20802
rect 19122 20750 19124 20802
rect 18844 20692 18900 20702
rect 18844 20598 18900 20636
rect 19068 20692 19124 20750
rect 18844 20244 18900 20254
rect 19068 20244 19124 20636
rect 18844 20242 19124 20244
rect 18844 20190 18846 20242
rect 18898 20190 19124 20242
rect 18844 20188 19124 20190
rect 18844 20178 18900 20188
rect 18508 20132 18564 20142
rect 18508 20130 18788 20132
rect 18508 20078 18510 20130
rect 18562 20078 18788 20130
rect 18508 20076 18788 20078
rect 18508 20066 18564 20076
rect 17052 19394 17108 19404
rect 18620 19346 18676 19358
rect 18620 19294 18622 19346
rect 18674 19294 18676 19346
rect 18508 18564 18564 18574
rect 18620 18564 18676 19294
rect 18508 18562 18676 18564
rect 18508 18510 18510 18562
rect 18562 18510 18676 18562
rect 18508 18508 18676 18510
rect 18508 18498 18564 18508
rect 18396 18228 18452 18238
rect 15820 16884 15876 16894
rect 15820 16790 15876 16828
rect 16604 16884 16660 16894
rect 16716 16884 16772 16940
rect 17724 18226 18452 18228
rect 17724 18174 18398 18226
rect 18450 18174 18452 18226
rect 17724 18172 18452 18174
rect 16604 16882 16772 16884
rect 16604 16830 16606 16882
rect 16658 16830 16772 16882
rect 16604 16828 16772 16830
rect 17388 16884 17444 16894
rect 16604 16818 16660 16828
rect 17388 16790 17444 16828
rect 17724 16882 17780 18172
rect 18396 18162 18452 18172
rect 18172 17108 18228 17118
rect 18732 17108 18788 20076
rect 18172 17014 18228 17052
rect 18284 17052 19012 17108
rect 17724 16830 17726 16882
rect 17778 16830 17780 16882
rect 16380 16658 16436 16670
rect 16380 16606 16382 16658
rect 16434 16606 16436 16658
rect 16268 16100 16324 16110
rect 16268 16006 16324 16044
rect 15372 15986 15540 15988
rect 15372 15934 15374 15986
rect 15426 15934 15540 15986
rect 15372 15932 15540 15934
rect 15596 15988 15652 15998
rect 15372 15922 15428 15932
rect 15596 15894 15652 15932
rect 16380 15876 16436 16606
rect 16492 16324 16548 16334
rect 16492 16230 16548 16268
rect 16716 16212 16772 16222
rect 16716 16098 16772 16156
rect 16716 16046 16718 16098
rect 16770 16046 16772 16098
rect 16716 16034 16772 16046
rect 17500 16100 17556 16110
rect 17500 16006 17556 16044
rect 17724 16098 17780 16830
rect 18060 16884 18116 16894
rect 17836 16660 17892 16670
rect 17836 16566 17892 16604
rect 17724 16046 17726 16098
rect 17778 16046 17780 16098
rect 17724 16034 17780 16046
rect 16940 15986 16996 15998
rect 16940 15934 16942 15986
rect 16994 15934 16996 15986
rect 16492 15876 16548 15886
rect 16380 15874 16548 15876
rect 16380 15822 16494 15874
rect 16546 15822 16548 15874
rect 16380 15820 16548 15822
rect 15148 15202 15204 15820
rect 16492 15810 16548 15820
rect 15148 15150 15150 15202
rect 15202 15150 15204 15202
rect 15148 15148 15204 15150
rect 16492 15204 16548 15242
rect 15148 15092 15428 15148
rect 16492 15092 16548 15148
rect 15036 14642 15092 14654
rect 15036 14590 15038 14642
rect 15090 14590 15092 14642
rect 14476 13346 14532 13356
rect 14812 13412 14868 13422
rect 14364 13134 14366 13186
rect 14418 13134 14420 13186
rect 14364 13122 14420 13134
rect 13916 12964 13972 12974
rect 13916 12870 13972 12908
rect 14252 12964 14308 12974
rect 14252 12870 14308 12908
rect 14476 12962 14532 12974
rect 14476 12910 14478 12962
rect 14530 12910 14532 12962
rect 14476 12516 14532 12910
rect 14028 12460 14532 12516
rect 14700 12738 14756 12750
rect 14700 12686 14702 12738
rect 14754 12686 14756 12738
rect 14028 12402 14084 12460
rect 14028 12350 14030 12402
rect 14082 12350 14084 12402
rect 14028 12338 14084 12350
rect 13916 12290 13972 12302
rect 13916 12238 13918 12290
rect 13970 12238 13972 12290
rect 12460 12180 12516 12190
rect 12460 12086 12516 12124
rect 12908 12178 12964 12190
rect 12908 12126 12910 12178
rect 12962 12126 12964 12178
rect 12908 12068 12964 12126
rect 13468 12180 13524 12190
rect 13468 12086 13524 12124
rect 12908 12002 12964 12012
rect 12572 11956 12628 11966
rect 12348 11900 12572 11956
rect 12572 11862 12628 11900
rect 13356 11732 13412 11742
rect 12796 11284 12852 11294
rect 12796 10722 12852 11228
rect 13244 10836 13300 10846
rect 13244 10742 13300 10780
rect 12796 10670 12798 10722
rect 12850 10670 12852 10722
rect 12796 10658 12852 10670
rect 12572 10612 12628 10622
rect 12572 10518 12628 10556
rect 12236 10334 12238 10386
rect 12290 10334 12292 10386
rect 12236 10322 12292 10334
rect 13356 10500 13412 11676
rect 12012 9938 12180 9940
rect 12012 9886 12014 9938
rect 12066 9886 12180 9938
rect 12012 9884 12180 9886
rect 12012 9874 12068 9884
rect 10668 9102 10670 9154
rect 10722 9102 10724 9154
rect 10668 9090 10724 9102
rect 11340 9268 11396 9278
rect 9884 8990 9886 9042
rect 9938 8990 9940 9042
rect 9884 8978 9940 8990
rect 11340 8484 11396 9212
rect 13244 9268 13300 9278
rect 13356 9268 13412 10444
rect 13916 10612 13972 12238
rect 14140 12292 14196 12302
rect 14140 12198 14196 12236
rect 14588 12290 14644 12302
rect 14588 12238 14590 12290
rect 14642 12238 14644 12290
rect 14476 12068 14532 12078
rect 14476 11974 14532 12012
rect 14588 11732 14644 12238
rect 14588 11666 14644 11676
rect 14364 11620 14420 11630
rect 14364 11394 14420 11564
rect 14476 11508 14532 11518
rect 14700 11508 14756 12686
rect 14812 12292 14868 13356
rect 14812 12198 14868 12236
rect 14476 11506 14756 11508
rect 14476 11454 14478 11506
rect 14530 11454 14756 11506
rect 14476 11452 14756 11454
rect 15036 11508 15092 14590
rect 15148 12964 15204 12974
rect 15148 12870 15204 12908
rect 15260 11956 15316 11966
rect 15148 11508 15204 11518
rect 15036 11452 15148 11508
rect 14476 11442 14532 11452
rect 15148 11442 15204 11452
rect 14364 11342 14366 11394
rect 14418 11342 14420 11394
rect 14364 11330 14420 11342
rect 14812 11396 14868 11406
rect 15260 11396 15316 11900
rect 15372 11508 15428 15092
rect 16268 15036 16492 15092
rect 16268 14530 16324 15036
rect 16492 15026 16548 15036
rect 16828 15092 16884 15102
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 16268 14466 16324 14478
rect 16604 14980 16660 14990
rect 16604 14532 16660 14924
rect 16604 14438 16660 14476
rect 15596 13970 15652 13982
rect 15596 13918 15598 13970
rect 15650 13918 15652 13970
rect 15484 13412 15540 13422
rect 15484 13186 15540 13356
rect 15484 13134 15486 13186
rect 15538 13134 15540 13186
rect 15484 13122 15540 13134
rect 15596 11618 15652 13918
rect 16156 13972 16212 13982
rect 16828 13972 16884 15036
rect 16940 14532 16996 15934
rect 17052 15988 17108 15998
rect 17052 15148 17108 15932
rect 17388 15988 17444 15998
rect 17388 15894 17444 15932
rect 17052 15092 17220 15148
rect 16940 14476 17108 14532
rect 16940 14308 16996 14318
rect 16940 14214 16996 14252
rect 16940 13972 16996 13982
rect 16828 13970 16996 13972
rect 16828 13918 16942 13970
rect 16994 13918 16996 13970
rect 16828 13916 16996 13918
rect 16156 13858 16212 13916
rect 16940 13906 16996 13916
rect 16156 13806 16158 13858
rect 16210 13806 16212 13858
rect 16156 13794 16212 13806
rect 16380 13860 16436 13870
rect 16380 13766 16436 13804
rect 17052 13860 17108 14476
rect 17164 14308 17220 15092
rect 17276 14532 17332 14542
rect 17276 14438 17332 14476
rect 17164 14242 17220 14252
rect 17612 14306 17668 14318
rect 17612 14254 17614 14306
rect 17666 14254 17668 14306
rect 17052 13794 17108 13804
rect 17612 13860 17668 14254
rect 17612 13794 17668 13804
rect 17724 13972 17780 13982
rect 15820 13746 15876 13758
rect 15820 13694 15822 13746
rect 15874 13694 15876 13746
rect 15820 13186 15876 13694
rect 15932 13748 15988 13758
rect 15932 13654 15988 13692
rect 17612 13636 17668 13646
rect 17724 13636 17780 13916
rect 17612 13634 17780 13636
rect 17612 13582 17614 13634
rect 17666 13582 17780 13634
rect 17612 13580 17780 13582
rect 17612 13570 17668 13580
rect 15820 13134 15822 13186
rect 15874 13134 15876 13186
rect 15820 13122 15876 13134
rect 15820 12964 15876 12974
rect 15820 12962 15988 12964
rect 15820 12910 15822 12962
rect 15874 12910 15988 12962
rect 15820 12908 15988 12910
rect 15820 12898 15876 12908
rect 15596 11566 15598 11618
rect 15650 11566 15652 11618
rect 15596 11554 15652 11566
rect 15932 11620 15988 12908
rect 18060 12962 18116 16828
rect 18172 16884 18228 16894
rect 18284 16884 18340 17052
rect 18172 16882 18340 16884
rect 18172 16830 18174 16882
rect 18226 16830 18340 16882
rect 18172 16828 18340 16830
rect 18620 16882 18676 16894
rect 18620 16830 18622 16882
rect 18674 16830 18676 16882
rect 18172 16818 18228 16828
rect 18620 16772 18676 16830
rect 18620 16706 18676 16716
rect 18508 16660 18564 16670
rect 18172 16212 18228 16222
rect 18172 16118 18228 16156
rect 18508 15538 18564 16604
rect 18508 15486 18510 15538
rect 18562 15486 18564 15538
rect 18508 15474 18564 15486
rect 18620 15428 18676 15438
rect 18620 15334 18676 15372
rect 18396 15314 18452 15326
rect 18396 15262 18398 15314
rect 18450 15262 18452 15314
rect 18396 15148 18452 15262
rect 18284 15092 18452 15148
rect 18844 15204 18900 15242
rect 18844 15138 18900 15148
rect 18284 13860 18340 15092
rect 18284 13766 18340 13804
rect 18396 14532 18452 14542
rect 18060 12910 18062 12962
rect 18114 12910 18116 12962
rect 18060 12898 18116 12910
rect 18396 12962 18452 14476
rect 18732 14420 18788 14430
rect 18732 14418 18900 14420
rect 18732 14366 18734 14418
rect 18786 14366 18900 14418
rect 18732 14364 18900 14366
rect 18732 14354 18788 14364
rect 18844 14308 18900 14364
rect 18620 13970 18676 13982
rect 18620 13918 18622 13970
rect 18674 13918 18676 13970
rect 18508 13748 18564 13758
rect 18508 13654 18564 13692
rect 18620 13186 18676 13918
rect 18732 13636 18788 13646
rect 18732 13542 18788 13580
rect 18844 13524 18900 14252
rect 18844 13458 18900 13468
rect 18620 13134 18622 13186
rect 18674 13134 18676 13186
rect 18620 13122 18676 13134
rect 18396 12910 18398 12962
rect 18450 12910 18452 12962
rect 18396 12898 18452 12910
rect 18844 12964 18900 12974
rect 18956 12964 19012 17052
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 19068 14754 19124 15262
rect 19068 14702 19070 14754
rect 19122 14702 19124 14754
rect 19068 14690 19124 14702
rect 19068 14532 19124 14542
rect 19068 14438 19124 14476
rect 19068 13746 19124 13758
rect 19068 13694 19070 13746
rect 19122 13694 19124 13746
rect 19068 13636 19124 13694
rect 19068 13570 19124 13580
rect 18844 12962 19012 12964
rect 18844 12910 18846 12962
rect 18898 12910 19012 12962
rect 18844 12908 19012 12910
rect 18172 12740 18228 12750
rect 15372 11452 15540 11508
rect 15260 11340 15428 11396
rect 14812 11302 14868 11340
rect 14028 11284 14084 11294
rect 14028 11190 14084 11228
rect 15148 11284 15204 11294
rect 15148 11190 15204 11228
rect 15372 11282 15428 11340
rect 15372 11230 15374 11282
rect 15426 11230 15428 11282
rect 15372 11218 15428 11230
rect 13244 9266 13412 9268
rect 13244 9214 13246 9266
rect 13298 9214 13412 9266
rect 13244 9212 13412 9214
rect 13692 9604 13748 9614
rect 13244 9202 13300 9212
rect 13692 9042 13748 9548
rect 13692 8990 13694 9042
rect 13746 8990 13748 9042
rect 13692 8978 13748 8990
rect 12796 8932 12852 8942
rect 13132 8932 13188 8942
rect 12796 8930 13188 8932
rect 12796 8878 12798 8930
rect 12850 8878 13134 8930
rect 13186 8878 13188 8930
rect 12796 8876 13188 8878
rect 12796 8866 12852 8876
rect 13132 8866 13188 8876
rect 9548 8036 9604 8046
rect 9548 7942 9604 7980
rect 10780 8036 10836 8046
rect 9044 7644 9156 7700
rect 8988 7606 9044 7644
rect 8204 7588 8260 7598
rect 7980 7586 8260 7588
rect 7980 7534 8206 7586
rect 8258 7534 8260 7586
rect 7980 7532 8260 7534
rect 8204 7522 8260 7532
rect 8540 7474 8596 7486
rect 8540 7422 8542 7474
rect 8594 7422 8596 7474
rect 8540 6802 8596 7422
rect 8540 6750 8542 6802
rect 8594 6750 8596 6802
rect 8540 6738 8596 6750
rect 7756 6638 7758 6690
rect 7810 6638 7812 6690
rect 7756 6626 7812 6638
rect 10780 6466 10836 7980
rect 10780 6414 10782 6466
rect 10834 6414 10836 6466
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 3612 4228 3668 4238
rect 3276 4226 3668 4228
rect 3276 4174 3614 4226
rect 3666 4174 3668 4226
rect 3276 4172 3668 4174
rect 2716 3444 2772 3454
rect 2940 3444 2996 3454
rect 2716 3442 2996 3444
rect 2716 3390 2718 3442
rect 2770 3390 2942 3442
rect 2994 3390 2996 3442
rect 2716 3388 2996 3390
rect 2716 800 2772 3388
rect 2940 3378 2996 3388
rect 3276 3442 3332 4172
rect 3612 4162 3668 4172
rect 3724 4228 3780 4238
rect 3724 4134 3780 4172
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 10780 3556 10836 6414
rect 11340 6690 11396 8428
rect 13356 8484 13412 8494
rect 13356 8372 13636 8428
rect 13580 8370 13636 8372
rect 13580 8318 13582 8370
rect 13634 8318 13636 8370
rect 11340 6638 11342 6690
rect 11394 6638 11396 6690
rect 11340 5906 11396 6638
rect 12124 7588 12180 7598
rect 12124 6018 12180 7532
rect 13580 6692 13636 8318
rect 13916 7698 13972 10556
rect 13916 7646 13918 7698
rect 13970 7646 13972 7698
rect 13916 7634 13972 7646
rect 14140 11170 14196 11182
rect 14140 11118 14142 11170
rect 14194 11118 14196 11170
rect 14140 7588 14196 11118
rect 14364 11172 14420 11182
rect 14364 9154 14420 11116
rect 15260 11172 15316 11182
rect 15260 11078 15316 11116
rect 15484 9604 15540 11452
rect 15820 11396 15876 11406
rect 15820 11302 15876 11340
rect 15932 10050 15988 11564
rect 17724 12738 18228 12740
rect 17724 12686 18174 12738
rect 18226 12686 18228 12738
rect 17724 12684 18228 12686
rect 16604 11508 16660 11518
rect 16604 11172 16660 11452
rect 17724 11506 17780 12684
rect 18172 12674 18228 12684
rect 17724 11454 17726 11506
rect 17778 11454 17780 11506
rect 17724 11442 17780 11454
rect 16940 11394 16996 11406
rect 16940 11342 16942 11394
rect 16994 11342 16996 11394
rect 16940 11172 16996 11342
rect 18844 11396 18900 12908
rect 19180 12404 19236 21420
rect 19292 17108 19348 17118
rect 19292 16994 19348 17052
rect 19292 16942 19294 16994
rect 19346 16942 19348 16994
rect 19292 16930 19348 16942
rect 19292 15428 19348 15438
rect 19404 15428 19460 25116
rect 19516 24834 19572 25230
rect 19740 25284 19796 25322
rect 19740 25218 19796 25228
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 19516 24782 19518 24834
rect 19570 24782 19572 24834
rect 19516 24770 19572 24782
rect 19740 24946 19796 24958
rect 19740 24894 19742 24946
rect 19794 24894 19796 24946
rect 19740 24052 19796 24894
rect 19852 24724 19908 24734
rect 19852 24630 19908 24668
rect 20076 24724 20132 24734
rect 20188 24724 20244 27022
rect 20300 29540 20356 29550
rect 20300 28642 20356 29484
rect 20412 29538 20468 29932
rect 20412 29486 20414 29538
rect 20466 29486 20468 29538
rect 20412 29474 20468 29486
rect 20300 28590 20302 28642
rect 20354 28590 20356 28642
rect 20300 26964 20356 28590
rect 20412 29092 20468 29102
rect 20412 28530 20468 29036
rect 20412 28478 20414 28530
rect 20466 28478 20468 28530
rect 20412 28466 20468 28478
rect 20524 28084 20580 30158
rect 20860 30212 20916 30222
rect 21196 30212 21252 30222
rect 20860 30210 21252 30212
rect 20860 30158 20862 30210
rect 20914 30158 21198 30210
rect 21250 30158 21252 30210
rect 20860 30156 21252 30158
rect 20860 30146 20916 30156
rect 21196 30146 21252 30156
rect 21532 30210 21588 30222
rect 21532 30158 21534 30210
rect 21586 30158 21588 30210
rect 20636 30100 20692 30110
rect 20636 30006 20692 30044
rect 21420 29988 21476 29998
rect 21420 29894 21476 29932
rect 21532 29316 21588 30158
rect 20636 29260 21588 29316
rect 20636 28642 20692 29260
rect 21420 29092 21476 29102
rect 21420 28754 21476 29036
rect 21420 28702 21422 28754
rect 21474 28702 21476 28754
rect 21420 28690 21476 28702
rect 20636 28590 20638 28642
rect 20690 28590 20692 28642
rect 20636 28578 20692 28590
rect 20524 28018 20580 28028
rect 20356 26908 20692 26964
rect 20300 26898 20356 26908
rect 20300 25284 20356 25294
rect 20300 25190 20356 25228
rect 20524 25172 20580 25182
rect 20524 24946 20580 25116
rect 20524 24894 20526 24946
rect 20578 24894 20580 24946
rect 20076 24722 20244 24724
rect 20076 24670 20078 24722
rect 20130 24670 20244 24722
rect 20076 24668 20244 24670
rect 20300 24724 20356 24734
rect 19964 24052 20020 24062
rect 19740 24050 20020 24052
rect 19740 23998 19966 24050
rect 20018 23998 20020 24050
rect 19740 23996 20020 23998
rect 19964 23986 20020 23996
rect 20076 23716 20132 24668
rect 20300 24630 20356 24668
rect 20076 23650 20132 23660
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 20412 22148 20468 22158
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 19628 21588 19684 21598
rect 20076 21588 20132 21598
rect 19628 21586 20132 21588
rect 19628 21534 19630 21586
rect 19682 21534 20078 21586
rect 20130 21534 20132 21586
rect 19628 21532 20132 21534
rect 19628 20692 19684 21532
rect 20076 21522 20132 21532
rect 20412 20916 20468 22092
rect 19964 20914 20468 20916
rect 19964 20862 20414 20914
rect 20466 20862 20468 20914
rect 19964 20860 20468 20862
rect 19964 20802 20020 20860
rect 20412 20850 20468 20860
rect 19964 20750 19966 20802
rect 20018 20750 20020 20802
rect 19964 20738 20020 20750
rect 19628 20598 19684 20636
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19852 18452 19908 18462
rect 19628 18450 19908 18452
rect 19628 18398 19854 18450
rect 19906 18398 19908 18450
rect 19628 18396 19908 18398
rect 19628 16772 19684 18396
rect 19852 18386 19908 18396
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19628 16706 19684 16716
rect 20524 16212 20580 24894
rect 20636 24836 20692 26908
rect 21644 26908 21700 32284
rect 21868 30212 21924 33182
rect 21868 30118 21924 30156
rect 21980 30884 22036 30894
rect 21756 28756 21812 28766
rect 21756 28084 21812 28700
rect 21980 28420 22036 30828
rect 21980 28354 22036 28364
rect 21868 28084 21924 28094
rect 21756 28082 22036 28084
rect 21756 28030 21870 28082
rect 21922 28030 22036 28082
rect 21756 28028 22036 28030
rect 21868 28018 21924 28028
rect 21980 27972 22036 28028
rect 21644 26852 21812 26908
rect 21084 25172 21140 25182
rect 21084 24946 21140 25116
rect 21084 24894 21086 24946
rect 21138 24894 21140 24946
rect 21084 24882 21140 24894
rect 20636 24742 20692 24780
rect 20748 23940 20804 23950
rect 21644 23940 21700 23950
rect 20748 23938 21700 23940
rect 20748 23886 20750 23938
rect 20802 23886 21646 23938
rect 21698 23886 21700 23938
rect 20748 23884 21700 23886
rect 20636 23492 20692 23502
rect 20636 22932 20692 23436
rect 20748 23044 20804 23884
rect 21644 23874 21700 23884
rect 21420 23716 21476 23726
rect 20972 23044 21028 23054
rect 20748 23042 21028 23044
rect 20748 22990 20974 23042
rect 21026 22990 21028 23042
rect 20748 22988 21028 22990
rect 20636 21586 20692 22876
rect 20636 21534 20638 21586
rect 20690 21534 20692 21586
rect 20636 21522 20692 21534
rect 20972 20244 21028 22988
rect 21420 22258 21476 23660
rect 21756 22372 21812 26852
rect 21980 26514 22036 27916
rect 21980 26462 21982 26514
rect 22034 26462 22036 26514
rect 21980 26450 22036 26462
rect 21868 24948 21924 24958
rect 21868 24854 21924 24892
rect 22092 23492 22148 40684
rect 22652 40740 22708 40750
rect 22316 40628 22372 40638
rect 22316 38946 22372 40572
rect 22652 40626 22708 40684
rect 22652 40574 22654 40626
rect 22706 40574 22708 40626
rect 22652 40562 22708 40574
rect 22316 38894 22318 38946
rect 22370 38894 22372 38946
rect 22316 38882 22372 38894
rect 22876 36932 22932 43820
rect 22988 41972 23044 41982
rect 22988 41300 23044 41916
rect 23324 41970 23380 44044
rect 23436 44034 23492 44044
rect 23660 42866 23716 42878
rect 23660 42814 23662 42866
rect 23714 42814 23716 42866
rect 23548 42530 23604 42542
rect 23548 42478 23550 42530
rect 23602 42478 23604 42530
rect 23548 42420 23604 42478
rect 23324 41918 23326 41970
rect 23378 41918 23380 41970
rect 23324 41906 23380 41918
rect 23436 42364 23604 42420
rect 23436 41972 23492 42364
rect 23436 41906 23492 41916
rect 23548 42196 23604 42206
rect 23660 42196 23716 42814
rect 24108 42754 24164 42766
rect 24108 42702 24110 42754
rect 24162 42702 24164 42754
rect 23772 42530 23828 42542
rect 23772 42478 23774 42530
rect 23826 42478 23828 42530
rect 23772 42420 23828 42478
rect 23772 42364 24052 42420
rect 23548 42194 23716 42196
rect 23548 42142 23550 42194
rect 23602 42142 23716 42194
rect 23548 42140 23716 42142
rect 22988 41234 23044 41244
rect 23100 41746 23156 41758
rect 23100 41694 23102 41746
rect 23154 41694 23156 41746
rect 22988 40516 23044 40526
rect 23100 40516 23156 41694
rect 23436 41748 23492 41758
rect 23436 41074 23492 41692
rect 23436 41022 23438 41074
rect 23490 41022 23492 41074
rect 23436 41010 23492 41022
rect 23436 40740 23492 40750
rect 23324 40628 23380 40638
rect 23324 40534 23380 40572
rect 22988 40514 23156 40516
rect 22988 40462 22990 40514
rect 23042 40462 23156 40514
rect 22988 40460 23156 40462
rect 22988 40450 23044 40460
rect 23324 40404 23380 40414
rect 23324 40310 23380 40348
rect 23436 40402 23492 40684
rect 23436 40350 23438 40402
rect 23490 40350 23492 40402
rect 23436 40338 23492 40350
rect 23548 40404 23604 42140
rect 23884 42084 23940 42094
rect 23772 41972 23828 41982
rect 23772 41878 23828 41916
rect 23884 41970 23940 42028
rect 23884 41918 23886 41970
rect 23938 41918 23940 41970
rect 23884 41906 23940 41918
rect 23660 41858 23716 41870
rect 23660 41806 23662 41858
rect 23714 41806 23716 41858
rect 23660 41188 23716 41806
rect 23660 41122 23716 41132
rect 23996 41524 24052 42364
rect 24108 42084 24164 42702
rect 24108 42028 24724 42084
rect 24444 41860 24500 41870
rect 24668 41860 24724 42028
rect 24444 41858 24612 41860
rect 24444 41806 24446 41858
rect 24498 41806 24612 41858
rect 24444 41804 24612 41806
rect 24444 41794 24500 41804
rect 24332 41748 24388 41758
rect 23996 40964 24052 41468
rect 23996 40898 24052 40908
rect 24108 41746 24388 41748
rect 24108 41694 24334 41746
rect 24386 41694 24388 41746
rect 24108 41692 24388 41694
rect 24108 40740 24164 41692
rect 24332 41682 24388 41692
rect 23884 40684 24164 40740
rect 24220 41300 24276 41310
rect 23884 40514 23940 40684
rect 24220 40516 24276 41244
rect 24556 41074 24612 41804
rect 24668 41794 24724 41804
rect 24780 41298 24836 45500
rect 24780 41246 24782 41298
rect 24834 41246 24836 41298
rect 24780 41234 24836 41246
rect 24556 41022 24558 41074
rect 24610 41022 24612 41074
rect 24332 40628 24388 40638
rect 24556 40628 24612 41022
rect 24332 40626 24612 40628
rect 24332 40574 24334 40626
rect 24386 40574 24612 40626
rect 24332 40572 24612 40574
rect 24332 40562 24388 40572
rect 23884 40462 23886 40514
rect 23938 40462 23940 40514
rect 23884 40450 23940 40462
rect 23996 40514 24276 40516
rect 23996 40462 24222 40514
rect 24274 40462 24276 40514
rect 23996 40460 24276 40462
rect 23660 40404 23716 40414
rect 23548 40402 23716 40404
rect 23548 40350 23662 40402
rect 23714 40350 23716 40402
rect 23548 40348 23716 40350
rect 23660 40338 23716 40348
rect 23996 39730 24052 40460
rect 24220 40450 24276 40460
rect 23996 39678 23998 39730
rect 24050 39678 24052 39730
rect 23996 39666 24052 39678
rect 24444 38722 24500 40572
rect 24556 40404 24612 40414
rect 24556 40310 24612 40348
rect 24444 38670 24446 38722
rect 24498 38670 24500 38722
rect 24444 38052 24500 38670
rect 24892 38668 24948 47292
rect 25004 48580 25060 48590
rect 25004 47460 25060 48524
rect 25228 48244 25284 48254
rect 25228 48150 25284 48188
rect 25340 47796 25396 48972
rect 25676 48692 25732 49758
rect 25676 48626 25732 48636
rect 25788 49810 25844 50372
rect 25788 49758 25790 49810
rect 25842 49758 25844 49810
rect 25676 48468 25732 48478
rect 25788 48468 25844 49758
rect 26460 49812 26516 49822
rect 26460 49810 26628 49812
rect 26460 49758 26462 49810
rect 26514 49758 26628 49810
rect 26460 49756 26628 49758
rect 26460 49746 26516 49756
rect 25676 48466 25844 48468
rect 25676 48414 25678 48466
rect 25730 48414 25844 48466
rect 25676 48412 25844 48414
rect 26572 48468 26628 49756
rect 26684 49810 26740 49822
rect 26684 49758 26686 49810
rect 26738 49758 26740 49810
rect 26684 49028 26740 49758
rect 26796 49698 26852 50540
rect 27132 50530 27188 50540
rect 27692 50596 27748 50606
rect 27356 50484 27412 50494
rect 27356 50390 27412 50428
rect 27580 50482 27636 50494
rect 27580 50430 27582 50482
rect 27634 50430 27636 50482
rect 27580 50034 27636 50430
rect 27580 49982 27582 50034
rect 27634 49982 27636 50034
rect 27580 49970 27636 49982
rect 26796 49646 26798 49698
rect 26850 49646 26852 49698
rect 26796 49634 26852 49646
rect 26908 49922 26964 49934
rect 26908 49870 26910 49922
rect 26962 49870 26964 49922
rect 26908 49476 26964 49870
rect 27356 49922 27412 49934
rect 27356 49870 27358 49922
rect 27410 49870 27412 49922
rect 26796 49420 26964 49476
rect 27244 49810 27300 49822
rect 27244 49758 27246 49810
rect 27298 49758 27300 49810
rect 26796 49252 26852 49420
rect 27244 49364 27300 49758
rect 27244 49298 27300 49308
rect 27356 49476 27412 49870
rect 27132 49252 27188 49262
rect 26796 49250 27188 49252
rect 26796 49198 27134 49250
rect 27186 49198 27188 49250
rect 26796 49196 27188 49198
rect 27132 49186 27188 49196
rect 27244 49140 27300 49150
rect 27356 49140 27412 49420
rect 27244 49138 27412 49140
rect 27244 49086 27246 49138
rect 27298 49086 27412 49138
rect 27244 49084 27412 49086
rect 27244 49074 27300 49084
rect 26684 48962 26740 48972
rect 27020 49028 27076 49038
rect 25676 48402 25732 48412
rect 25564 48356 25620 48366
rect 25564 48262 25620 48300
rect 25228 47740 25396 47796
rect 25788 48242 25844 48254
rect 25788 48190 25790 48242
rect 25842 48190 25844 48242
rect 25116 47460 25172 47470
rect 25004 47458 25172 47460
rect 25004 47406 25118 47458
rect 25170 47406 25172 47458
rect 25004 47404 25172 47406
rect 25004 45778 25060 47404
rect 25116 47394 25172 47404
rect 25004 45726 25006 45778
rect 25058 45726 25060 45778
rect 25004 45714 25060 45726
rect 25228 45332 25284 47740
rect 25340 47572 25396 47582
rect 25788 47572 25844 48190
rect 26236 48244 26292 48254
rect 26460 48244 26516 48254
rect 26292 48242 26516 48244
rect 26292 48190 26462 48242
rect 26514 48190 26516 48242
rect 26292 48188 26516 48190
rect 26236 48150 26292 48188
rect 26460 48178 26516 48188
rect 26572 47682 26628 48412
rect 27020 48916 27076 48972
rect 27020 48860 27412 48916
rect 27020 48466 27076 48860
rect 27132 48692 27188 48702
rect 27188 48636 27300 48692
rect 27132 48626 27188 48636
rect 27020 48414 27022 48466
rect 27074 48414 27076 48466
rect 27020 48402 27076 48414
rect 27132 48468 27188 48478
rect 27132 48374 27188 48412
rect 26572 47630 26574 47682
rect 26626 47630 26628 47682
rect 26012 47572 26068 47582
rect 25340 47570 25732 47572
rect 25340 47518 25342 47570
rect 25394 47518 25732 47570
rect 25340 47516 25732 47518
rect 25788 47516 26012 47572
rect 25340 47506 25396 47516
rect 25676 47458 25732 47516
rect 25676 47406 25678 47458
rect 25730 47406 25732 47458
rect 25676 47394 25732 47406
rect 26012 47458 26068 47516
rect 26012 47406 26014 47458
rect 26066 47406 26068 47458
rect 26012 47394 26068 47406
rect 26348 47460 26404 47470
rect 26348 47366 26404 47404
rect 25452 47348 25508 47358
rect 25452 47254 25508 47292
rect 26572 47348 26628 47630
rect 26572 47282 26628 47292
rect 26908 48356 26964 48366
rect 26908 48242 26964 48300
rect 27244 48244 27300 48636
rect 26908 48190 26910 48242
rect 26962 48190 26964 48242
rect 26236 47236 26292 47246
rect 26236 47142 26292 47180
rect 25452 45668 25508 45678
rect 25452 45574 25508 45612
rect 25228 44324 25284 45276
rect 26012 45108 26068 45118
rect 26012 45106 26516 45108
rect 26012 45054 26014 45106
rect 26066 45054 26516 45106
rect 26012 45052 26516 45054
rect 26012 45042 26068 45052
rect 26124 44884 26180 44894
rect 26124 44882 26404 44884
rect 26124 44830 26126 44882
rect 26178 44830 26404 44882
rect 26124 44828 26404 44830
rect 26124 44818 26180 44828
rect 25228 44258 25284 44268
rect 25452 44492 25956 44548
rect 25452 44322 25508 44492
rect 25900 44436 25956 44492
rect 26124 44436 26180 44446
rect 25900 44434 26180 44436
rect 25900 44382 26126 44434
rect 26178 44382 26180 44434
rect 25900 44380 26180 44382
rect 26124 44370 26180 44380
rect 25452 44270 25454 44322
rect 25506 44270 25508 44322
rect 25452 44258 25508 44270
rect 25564 44324 25620 44334
rect 25116 44210 25172 44222
rect 25116 44158 25118 44210
rect 25170 44158 25172 44210
rect 25116 43764 25172 44158
rect 25116 43698 25172 43708
rect 25452 44098 25508 44110
rect 25452 44046 25454 44098
rect 25506 44046 25508 44098
rect 25452 40516 25508 44046
rect 25564 43538 25620 44268
rect 25564 43486 25566 43538
rect 25618 43486 25620 43538
rect 25564 43474 25620 43486
rect 25788 44322 25844 44334
rect 25788 44270 25790 44322
rect 25842 44270 25844 44322
rect 25788 43426 25844 44270
rect 26012 44098 26068 44110
rect 26012 44046 26014 44098
rect 26066 44046 26068 44098
rect 25900 43540 25956 43550
rect 25900 43446 25956 43484
rect 25788 43374 25790 43426
rect 25842 43374 25844 43426
rect 25788 43362 25844 43374
rect 26012 43316 26068 44046
rect 26236 44100 26292 44110
rect 26236 44006 26292 44044
rect 26124 43764 26180 43774
rect 26348 43764 26404 44828
rect 26124 43762 26404 43764
rect 26124 43710 26126 43762
rect 26178 43710 26404 43762
rect 26124 43708 26404 43710
rect 26460 44098 26516 45052
rect 26908 44546 26964 48190
rect 27132 48188 27300 48244
rect 27020 47572 27076 47582
rect 27020 47458 27076 47516
rect 27020 47406 27022 47458
rect 27074 47406 27076 47458
rect 27020 47394 27076 47406
rect 27132 47458 27188 48188
rect 27132 47406 27134 47458
rect 27186 47406 27188 47458
rect 27132 47236 27188 47406
rect 27132 47170 27188 47180
rect 27244 47346 27300 47358
rect 27244 47294 27246 47346
rect 27298 47294 27300 47346
rect 27244 46900 27300 47294
rect 27244 46834 27300 46844
rect 27356 46786 27412 48860
rect 27580 48244 27636 48254
rect 27580 48150 27636 48188
rect 27692 47348 27748 50540
rect 28588 50484 28644 50494
rect 28588 49922 28644 50428
rect 28588 49870 28590 49922
rect 28642 49870 28644 49922
rect 28588 49858 28644 49870
rect 31052 49922 31108 49934
rect 31052 49870 31054 49922
rect 31106 49870 31108 49922
rect 27916 49810 27972 49822
rect 27916 49758 27918 49810
rect 27970 49758 27972 49810
rect 27916 48804 27972 49758
rect 30716 49698 30772 49710
rect 30716 49646 30718 49698
rect 30770 49646 30772 49698
rect 27916 48738 27972 48748
rect 28476 49476 28532 49486
rect 28252 47460 28308 47470
rect 28252 47366 28308 47404
rect 27916 47348 27972 47358
rect 27580 47346 27748 47348
rect 27580 47294 27694 47346
rect 27746 47294 27748 47346
rect 27580 47292 27748 47294
rect 27468 46900 27524 46910
rect 27468 46806 27524 46844
rect 27356 46734 27358 46786
rect 27410 46734 27412 46786
rect 27356 46722 27412 46734
rect 26908 44494 26910 44546
rect 26962 44494 26964 44546
rect 26908 44482 26964 44494
rect 26460 44046 26462 44098
rect 26514 44046 26516 44098
rect 26124 43698 26180 43708
rect 26012 43250 26068 43260
rect 26124 41972 26180 41982
rect 26012 41300 26068 41310
rect 26124 41300 26180 41916
rect 26348 41972 26404 41982
rect 26460 41972 26516 44046
rect 27020 44100 27076 44110
rect 27020 43708 27076 44044
rect 26796 43652 27076 43708
rect 27132 44098 27188 44110
rect 27132 44046 27134 44098
rect 27186 44046 27188 44098
rect 26796 43650 26852 43652
rect 26796 43598 26798 43650
rect 26850 43598 26852 43650
rect 26796 43586 26852 43598
rect 27132 43540 27188 44046
rect 27468 43764 27524 43774
rect 27580 43764 27636 47292
rect 27692 47282 27748 47292
rect 27804 47346 27972 47348
rect 27804 47294 27918 47346
rect 27970 47294 27972 47346
rect 27804 47292 27972 47294
rect 27692 46900 27748 46910
rect 27804 46900 27860 47292
rect 27916 47282 27972 47292
rect 28140 47348 28196 47358
rect 28140 47254 28196 47292
rect 27692 46898 27860 46900
rect 27692 46846 27694 46898
rect 27746 46846 27860 46898
rect 27692 46844 27860 46846
rect 27692 46834 27748 46844
rect 28476 46676 28532 49420
rect 30716 49476 30772 49646
rect 30716 49410 30772 49420
rect 27524 43708 27636 43764
rect 28364 44996 28420 45006
rect 28364 44660 28420 44940
rect 27468 43698 27524 43708
rect 27916 43652 27972 43662
rect 28364 43652 28420 44604
rect 27916 43650 28420 43652
rect 27916 43598 27918 43650
rect 27970 43598 28420 43650
rect 27916 43596 28420 43598
rect 27916 43586 27972 43596
rect 26908 43484 27132 43540
rect 26908 42196 26964 43484
rect 27132 43446 27188 43484
rect 27356 43538 27412 43550
rect 27356 43486 27358 43538
rect 27410 43486 27412 43538
rect 27244 43428 27300 43438
rect 27244 43334 27300 43372
rect 27356 43316 27412 43486
rect 28364 43538 28420 43596
rect 28364 43486 28366 43538
rect 28418 43486 28420 43538
rect 28364 43474 28420 43486
rect 28476 43316 28532 46620
rect 29148 48804 29204 48814
rect 29148 47458 29204 48748
rect 30940 48804 30996 48814
rect 30940 48710 30996 48748
rect 31052 48692 31108 49870
rect 31164 49812 31220 50652
rect 40348 50706 40404 50718
rect 40348 50654 40350 50706
rect 40402 50654 40404 50706
rect 33964 50596 34020 50606
rect 33964 50594 34132 50596
rect 33964 50542 33966 50594
rect 34018 50542 34132 50594
rect 33964 50540 34132 50542
rect 33964 50530 34020 50540
rect 33180 50484 33236 50494
rect 32060 50482 33236 50484
rect 32060 50430 33182 50482
rect 33234 50430 33236 50482
rect 32060 50428 33236 50430
rect 34076 50428 34132 50540
rect 37436 50594 37492 50606
rect 37436 50542 37438 50594
rect 37490 50542 37492 50594
rect 37436 50428 37492 50542
rect 31948 49922 32004 49934
rect 31948 49870 31950 49922
rect 32002 49870 32004 49922
rect 31276 49812 31332 49822
rect 31164 49810 31332 49812
rect 31164 49758 31278 49810
rect 31330 49758 31332 49810
rect 31164 49756 31332 49758
rect 31052 48626 31108 48636
rect 29148 47406 29150 47458
rect 29202 47406 29204 47458
rect 29148 44322 29204 47406
rect 29932 47348 29988 47358
rect 29932 47254 29988 47292
rect 31276 47124 31332 49756
rect 31724 49700 31780 49710
rect 31724 49606 31780 49644
rect 31948 49140 32004 49870
rect 32060 49698 32116 50428
rect 33180 50418 33236 50428
rect 32060 49646 32062 49698
rect 32114 49646 32116 49698
rect 32060 49634 32116 49646
rect 33964 50372 34468 50428
rect 33964 49810 34020 50372
rect 34412 50370 34468 50372
rect 34412 50318 34414 50370
rect 34466 50318 34468 50370
rect 34412 50306 34468 50318
rect 37100 50372 37492 50428
rect 38220 50484 38276 50494
rect 38220 50482 38500 50484
rect 38220 50430 38222 50482
rect 38274 50430 38500 50482
rect 38220 50428 38500 50430
rect 38220 50418 38276 50428
rect 37100 50370 37156 50372
rect 37100 50318 37102 50370
rect 37154 50318 37156 50370
rect 33964 49758 33966 49810
rect 34018 49758 34020 49810
rect 32060 49140 32116 49150
rect 31948 49084 32060 49140
rect 31948 48242 32004 49084
rect 32060 49074 32116 49084
rect 33964 48804 34020 49758
rect 34748 49700 34804 49710
rect 36876 49700 36932 49710
rect 34748 49698 35140 49700
rect 34748 49646 34750 49698
rect 34802 49646 35140 49698
rect 34748 49644 35140 49646
rect 34748 49634 34804 49644
rect 35084 49250 35140 49644
rect 36764 49698 36932 49700
rect 36764 49646 36878 49698
rect 36930 49646 36932 49698
rect 36764 49644 36932 49646
rect 35644 49476 35700 49486
rect 35196 49420 35460 49430
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35196 49354 35460 49364
rect 35532 49420 35644 49476
rect 35084 49198 35086 49250
rect 35138 49198 35140 49250
rect 35084 49186 35140 49198
rect 35420 49252 35476 49262
rect 35532 49252 35588 49420
rect 35644 49410 35700 49420
rect 35420 49250 35588 49252
rect 35420 49198 35422 49250
rect 35474 49198 35588 49250
rect 35420 49196 35588 49198
rect 35420 49186 35476 49196
rect 35196 49140 35252 49150
rect 35196 48914 35252 49084
rect 35196 48862 35198 48914
rect 35250 48862 35252 48914
rect 35196 48850 35252 48862
rect 36764 48916 36820 49644
rect 36876 49634 36932 49644
rect 36764 48850 36820 48860
rect 33964 48738 34020 48748
rect 35532 48804 35588 48814
rect 31948 48190 31950 48242
rect 32002 48190 32004 48242
rect 31948 48178 32004 48190
rect 32284 48692 32340 48702
rect 31612 48132 31668 48142
rect 31612 48038 31668 48076
rect 31948 48020 32004 48030
rect 31948 47926 32004 47964
rect 30828 47068 31332 47124
rect 32060 47570 32116 47582
rect 32060 47518 32062 47570
rect 32114 47518 32116 47570
rect 30268 46786 30324 46798
rect 30268 46734 30270 46786
rect 30322 46734 30324 46786
rect 30156 46674 30212 46686
rect 30156 46622 30158 46674
rect 30210 46622 30212 46674
rect 29932 46564 29988 46574
rect 29932 46470 29988 46508
rect 30156 46452 30212 46622
rect 30268 46676 30324 46734
rect 30268 46610 30324 46620
rect 30828 46452 30884 47068
rect 30156 46396 30884 46452
rect 30940 46900 30996 46910
rect 30940 46786 30996 46844
rect 32060 46900 32116 47518
rect 32060 46834 32116 46844
rect 32284 47460 32340 48636
rect 33180 48020 33236 48030
rect 33180 47570 33236 47964
rect 35196 47852 35460 47862
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35196 47786 35460 47796
rect 33180 47518 33182 47570
rect 33234 47518 33236 47570
rect 33180 47506 33236 47518
rect 33740 47572 33796 47582
rect 32396 47460 32452 47470
rect 32284 47458 32452 47460
rect 32284 47406 32398 47458
rect 32450 47406 32452 47458
rect 32284 47404 32452 47406
rect 32284 46900 32340 47404
rect 32396 47394 32452 47404
rect 32284 46898 32564 46900
rect 32284 46846 32286 46898
rect 32338 46846 32564 46898
rect 32284 46844 32564 46846
rect 32284 46834 32340 46844
rect 30940 46734 30942 46786
rect 30994 46734 30996 46786
rect 29148 44270 29150 44322
rect 29202 44270 29204 44322
rect 27356 43250 27412 43260
rect 28140 43260 28532 43316
rect 28588 43650 28644 43662
rect 28588 43598 28590 43650
rect 28642 43598 28644 43650
rect 28588 43540 28644 43598
rect 28588 43316 28644 43484
rect 27020 42196 27076 42206
rect 26348 41970 26516 41972
rect 26348 41918 26350 41970
rect 26402 41918 26516 41970
rect 26348 41916 26516 41918
rect 26796 42194 27076 42196
rect 26796 42142 27022 42194
rect 27074 42142 27076 42194
rect 26796 42140 27076 42142
rect 26796 41970 26852 42140
rect 27020 42130 27076 42140
rect 26796 41918 26798 41970
rect 26850 41918 26852 41970
rect 26348 41524 26404 41916
rect 26796 41906 26852 41918
rect 27356 41970 27412 41982
rect 27356 41918 27358 41970
rect 27410 41918 27412 41970
rect 26348 41458 26404 41468
rect 26572 41858 26628 41870
rect 26572 41806 26574 41858
rect 26626 41806 26628 41858
rect 26460 41412 26516 41422
rect 26572 41412 26628 41806
rect 27356 41860 27412 41918
rect 27356 41794 27412 41804
rect 26460 41410 26628 41412
rect 26460 41358 26462 41410
rect 26514 41358 26628 41410
rect 26460 41356 26628 41358
rect 26796 41412 26852 41422
rect 26460 41346 26516 41356
rect 26068 41244 26180 41300
rect 26012 41186 26068 41244
rect 26012 41134 26014 41186
rect 26066 41134 26068 41186
rect 26012 41122 26068 41134
rect 26572 41188 26628 41198
rect 26572 41094 26628 41132
rect 26460 40962 26516 40974
rect 26460 40910 26462 40962
rect 26514 40910 26516 40962
rect 26460 40516 26516 40910
rect 26796 40964 26852 41356
rect 27916 41300 27972 41310
rect 27356 40964 27412 40974
rect 26796 40962 27412 40964
rect 26796 40910 27358 40962
rect 27410 40910 27412 40962
rect 26796 40908 27412 40910
rect 26572 40516 26628 40526
rect 26460 40514 26628 40516
rect 26460 40462 26574 40514
rect 26626 40462 26628 40514
rect 26460 40460 26628 40462
rect 25452 40450 25508 40460
rect 26572 40450 26628 40460
rect 25900 40404 25956 40414
rect 25900 40310 25956 40348
rect 27356 38668 27412 40908
rect 27916 39730 27972 41244
rect 27916 39678 27918 39730
rect 27970 39678 27972 39730
rect 27916 39666 27972 39678
rect 24892 38612 25620 38668
rect 27356 38612 27524 38668
rect 24444 37986 24500 37996
rect 25340 37380 25396 37390
rect 25340 37156 25396 37324
rect 25564 37266 25620 38612
rect 25788 38052 25844 38062
rect 25788 37958 25844 37996
rect 26348 38052 26404 38062
rect 26348 37958 26404 37996
rect 26908 38052 26964 38062
rect 26460 37938 26516 37950
rect 26460 37886 26462 37938
rect 26514 37886 26516 37938
rect 26460 37604 26516 37886
rect 26460 37538 26516 37548
rect 26908 37826 26964 37996
rect 26908 37774 26910 37826
rect 26962 37774 26964 37826
rect 26796 37380 26852 37390
rect 26796 37286 26852 37324
rect 25564 37214 25566 37266
rect 25618 37214 25620 37266
rect 25564 37202 25620 37214
rect 26236 37268 26292 37278
rect 26236 37174 26292 37212
rect 22876 36866 22932 36876
rect 25228 37154 25396 37156
rect 25228 37102 25342 37154
rect 25394 37102 25396 37154
rect 25228 37100 25396 37102
rect 26908 37156 26964 37774
rect 26908 37100 27188 37156
rect 22316 36372 22372 36382
rect 22316 35922 22372 36316
rect 22428 36372 22484 36382
rect 24668 36372 24724 36382
rect 22428 36370 22932 36372
rect 22428 36318 22430 36370
rect 22482 36318 22932 36370
rect 22428 36316 22932 36318
rect 22428 36306 22484 36316
rect 22316 35870 22318 35922
rect 22370 35870 22372 35922
rect 22316 35858 22372 35870
rect 22876 35922 22932 36316
rect 24668 36258 24724 36316
rect 24668 36206 24670 36258
rect 24722 36206 24724 36258
rect 24668 36194 24724 36206
rect 22876 35870 22878 35922
rect 22930 35870 22932 35922
rect 22876 35858 22932 35870
rect 22540 35812 22596 35822
rect 22540 35810 22708 35812
rect 22540 35758 22542 35810
rect 22594 35758 22708 35810
rect 22540 35756 22708 35758
rect 22540 35746 22596 35756
rect 22204 35698 22260 35710
rect 22204 35646 22206 35698
rect 22258 35646 22260 35698
rect 22204 34916 22260 35646
rect 22652 35698 22708 35756
rect 22652 35646 22654 35698
rect 22706 35646 22708 35698
rect 22652 35634 22708 35646
rect 23100 35698 23156 35710
rect 23100 35646 23102 35698
rect 23154 35646 23156 35698
rect 22204 34850 22260 34860
rect 23100 33348 23156 35646
rect 23324 35698 23380 35710
rect 23324 35646 23326 35698
rect 23378 35646 23380 35698
rect 23324 35588 23380 35646
rect 23772 35588 23828 35598
rect 23324 35586 23828 35588
rect 23324 35534 23774 35586
rect 23826 35534 23828 35586
rect 23324 35532 23828 35534
rect 23772 34132 23828 35532
rect 24556 34916 24612 34926
rect 24556 34822 24612 34860
rect 24220 34692 24276 34702
rect 24220 34580 24276 34636
rect 24668 34690 24724 34702
rect 24668 34638 24670 34690
rect 24722 34638 24724 34690
rect 24668 34580 24724 34638
rect 24892 34692 24948 34702
rect 24892 34598 24948 34636
rect 24220 34524 24668 34580
rect 24668 34514 24724 34524
rect 23772 34066 23828 34076
rect 23324 34020 23380 34030
rect 23324 33926 23380 33964
rect 23996 34020 24052 34030
rect 23212 33348 23268 33358
rect 23100 33346 23268 33348
rect 23100 33294 23214 33346
rect 23266 33294 23268 33346
rect 23100 33292 23268 33294
rect 23212 33282 23268 33292
rect 22764 33236 22820 33246
rect 22764 32786 22820 33180
rect 23548 33236 23604 33246
rect 23548 33234 23716 33236
rect 23548 33182 23550 33234
rect 23602 33182 23716 33234
rect 23548 33180 23716 33182
rect 23548 33170 23604 33180
rect 23436 33124 23492 33134
rect 23436 33030 23492 33068
rect 23660 32788 23716 33180
rect 22764 32734 22766 32786
rect 22818 32734 22820 32786
rect 22764 32722 22820 32734
rect 23100 32732 23716 32788
rect 22988 32674 23044 32686
rect 22988 32622 22990 32674
rect 23042 32622 23044 32674
rect 22988 32564 23044 32622
rect 23100 32674 23156 32732
rect 23100 32622 23102 32674
rect 23154 32622 23156 32674
rect 23100 32610 23156 32622
rect 22988 32498 23044 32508
rect 23548 32564 23604 32574
rect 23548 32470 23604 32508
rect 23436 31892 23492 31902
rect 23436 31780 23492 31836
rect 23212 31778 23492 31780
rect 23212 31726 23438 31778
rect 23490 31726 23492 31778
rect 23212 31724 23492 31726
rect 22540 30100 22596 30110
rect 22428 29876 22484 29886
rect 22204 28084 22260 28094
rect 22204 27990 22260 28028
rect 22428 27636 22484 29820
rect 22540 29314 22596 30044
rect 23212 29652 23268 31724
rect 23436 31714 23492 31724
rect 23660 31668 23716 32732
rect 23996 31778 24052 33964
rect 24668 34020 24724 34030
rect 24780 34020 24836 34030
rect 24668 34018 24780 34020
rect 24668 33966 24670 34018
rect 24722 33966 24780 34018
rect 24668 33964 24780 33966
rect 24668 33954 24724 33964
rect 24108 33124 24164 33134
rect 24108 32676 24164 33068
rect 24108 32610 24164 32620
rect 24668 32450 24724 32462
rect 24668 32398 24670 32450
rect 24722 32398 24724 32450
rect 23996 31726 23998 31778
rect 24050 31726 24052 31778
rect 23996 31714 24052 31726
rect 24108 31836 24500 31892
rect 23660 31574 23716 31612
rect 23884 30436 23940 30446
rect 23884 30322 23940 30380
rect 23884 30270 23886 30322
rect 23938 30270 23940 30322
rect 23884 30258 23940 30270
rect 23996 30212 24052 30222
rect 24108 30212 24164 31836
rect 24444 31780 24500 31836
rect 24556 31780 24612 31790
rect 24444 31778 24612 31780
rect 24444 31726 24558 31778
rect 24610 31726 24612 31778
rect 24444 31724 24612 31726
rect 24556 31714 24612 31724
rect 24220 31554 24276 31566
rect 24220 31502 24222 31554
rect 24274 31502 24276 31554
rect 24220 31108 24276 31502
rect 24332 31554 24388 31566
rect 24332 31502 24334 31554
rect 24386 31502 24388 31554
rect 24332 31444 24388 31502
rect 24332 31378 24388 31388
rect 24444 31554 24500 31566
rect 24444 31502 24446 31554
rect 24498 31502 24500 31554
rect 24220 31042 24276 31052
rect 24444 31332 24500 31502
rect 24668 31332 24724 32398
rect 23996 30210 24164 30212
rect 23996 30158 23998 30210
rect 24050 30158 24164 30210
rect 23996 30156 24164 30158
rect 23324 30100 23380 30110
rect 23324 30006 23380 30044
rect 23212 29558 23268 29596
rect 23548 29986 23604 29998
rect 23772 29988 23828 29998
rect 23548 29934 23550 29986
rect 23602 29934 23604 29986
rect 22876 29540 22932 29550
rect 22876 29446 22932 29484
rect 22540 29262 22542 29314
rect 22594 29262 22596 29314
rect 22540 29250 22596 29262
rect 23436 28532 23492 28542
rect 22764 28028 23044 28084
rect 22428 27570 22484 27580
rect 22540 27858 22596 27870
rect 22540 27806 22542 27858
rect 22594 27806 22596 27858
rect 22204 27524 22260 27534
rect 22204 27076 22260 27468
rect 22540 27524 22596 27806
rect 22540 27458 22596 27468
rect 22204 24834 22260 27020
rect 22316 24948 22372 24958
rect 22316 24854 22372 24892
rect 22204 24782 22206 24834
rect 22258 24782 22260 24834
rect 22204 24770 22260 24782
rect 22652 24722 22708 24734
rect 22652 24670 22654 24722
rect 22706 24670 22708 24722
rect 22092 23426 22148 23436
rect 22316 24498 22372 24510
rect 22316 24446 22318 24498
rect 22370 24446 22372 24498
rect 22316 23154 22372 24446
rect 22428 23826 22484 23838
rect 22428 23774 22430 23826
rect 22482 23774 22484 23826
rect 22428 23380 22484 23774
rect 22540 23380 22596 23390
rect 22428 23378 22596 23380
rect 22428 23326 22542 23378
rect 22594 23326 22596 23378
rect 22428 23324 22596 23326
rect 22540 23314 22596 23324
rect 22316 23102 22318 23154
rect 22370 23102 22372 23154
rect 22316 23090 22372 23102
rect 22652 23154 22708 24670
rect 22652 23102 22654 23154
rect 22706 23102 22708 23154
rect 22652 23090 22708 23102
rect 21756 22306 21812 22316
rect 21420 22206 21422 22258
rect 21474 22206 21476 22258
rect 21420 22194 21476 22206
rect 21756 22146 21812 22158
rect 21756 22094 21758 22146
rect 21810 22094 21812 22146
rect 21756 21812 21812 22094
rect 21868 21812 21924 21822
rect 21756 21756 21868 21812
rect 21868 21718 21924 21756
rect 22204 21812 22260 21822
rect 21532 21586 21588 21598
rect 21532 21534 21534 21586
rect 21586 21534 21588 21586
rect 21532 21364 21588 21534
rect 21532 21298 21588 21308
rect 22204 20802 22260 21756
rect 22652 21812 22708 21822
rect 22652 21718 22708 21756
rect 22316 21474 22372 21486
rect 22316 21422 22318 21474
rect 22370 21422 22372 21474
rect 22316 21364 22372 21422
rect 22316 21298 22372 21308
rect 22204 20750 22206 20802
rect 22258 20750 22260 20802
rect 22204 20738 22260 20750
rect 20972 20178 21028 20188
rect 21868 20578 21924 20590
rect 21868 20526 21870 20578
rect 21922 20526 21924 20578
rect 21532 19012 21588 19022
rect 20636 18340 20692 18350
rect 20636 18338 21476 18340
rect 20636 18286 20638 18338
rect 20690 18286 21476 18338
rect 20636 18284 21476 18286
rect 20636 18274 20692 18284
rect 21420 17778 21476 18284
rect 21420 17726 21422 17778
rect 21474 17726 21476 17778
rect 21420 17714 21476 17726
rect 21308 17556 21364 17566
rect 21532 17556 21588 18956
rect 21868 17668 21924 20526
rect 22204 20244 22260 20254
rect 22092 19684 22148 19694
rect 22092 17780 22148 19628
rect 22092 17714 22148 17724
rect 22204 19012 22260 20188
rect 22764 19122 22820 28028
rect 22988 27970 23044 28028
rect 22988 27918 22990 27970
rect 23042 27918 23044 27970
rect 22988 27906 23044 27918
rect 23436 27860 23492 28476
rect 23436 27766 23492 27804
rect 23324 27076 23380 27086
rect 22988 27074 23380 27076
rect 22988 27022 23326 27074
rect 23378 27022 23380 27074
rect 22988 27020 23380 27022
rect 22988 26962 23044 27020
rect 23324 27010 23380 27020
rect 22988 26910 22990 26962
rect 23042 26910 23044 26962
rect 22988 25284 23044 26910
rect 23548 26962 23604 29934
rect 23548 26910 23550 26962
rect 23602 26910 23604 26962
rect 23548 26852 23604 26910
rect 23660 29932 23772 29988
rect 23660 26908 23716 29932
rect 23772 29894 23828 29932
rect 23996 28532 24052 30156
rect 23996 28466 24052 28476
rect 24332 28642 24388 28654
rect 24332 28590 24334 28642
rect 24386 28590 24388 28642
rect 23996 28084 24052 28094
rect 24220 28084 24276 28094
rect 24332 28084 24388 28590
rect 23996 27990 24052 28028
rect 24108 28082 24388 28084
rect 24108 28030 24222 28082
rect 24274 28030 24388 28082
rect 24108 28028 24388 28030
rect 23772 27972 23828 27982
rect 23772 27858 23828 27916
rect 23772 27806 23774 27858
rect 23826 27806 23828 27858
rect 23772 27794 23828 27806
rect 23660 26852 23828 26908
rect 23548 26786 23604 26796
rect 22988 25218 23044 25228
rect 22876 24834 22932 24846
rect 22876 24782 22878 24834
rect 22930 24782 22932 24834
rect 22876 24612 22932 24782
rect 22988 24836 23044 24846
rect 22988 24742 23044 24780
rect 23436 24612 23492 24622
rect 22876 24610 23492 24612
rect 22876 24558 23438 24610
rect 23490 24558 23492 24610
rect 22876 24556 23492 24558
rect 22988 23154 23044 23166
rect 22988 23102 22990 23154
rect 23042 23102 23044 23154
rect 22988 21700 23044 23102
rect 22988 21634 23044 21644
rect 23212 21588 23268 21598
rect 23212 21494 23268 21532
rect 23436 19684 23492 24556
rect 23660 22372 23716 22382
rect 23548 21812 23604 21822
rect 23548 21698 23604 21756
rect 23548 21646 23550 21698
rect 23602 21646 23604 21698
rect 23548 21634 23604 21646
rect 23660 20020 23716 22316
rect 23436 19618 23492 19628
rect 23548 19964 23716 20020
rect 23212 19234 23268 19246
rect 23212 19182 23214 19234
rect 23266 19182 23268 19234
rect 22764 19070 22766 19122
rect 22818 19070 22820 19122
rect 22316 19012 22372 19022
rect 22204 19010 22372 19012
rect 22204 18958 22318 19010
rect 22370 18958 22372 19010
rect 22204 18956 22372 18958
rect 21868 17574 21924 17612
rect 21308 17554 21588 17556
rect 21308 17502 21310 17554
rect 21362 17502 21588 17554
rect 21308 17500 21588 17502
rect 21644 17556 21700 17566
rect 21644 17554 21812 17556
rect 21644 17502 21646 17554
rect 21698 17502 21812 17554
rect 21644 17500 21812 17502
rect 21308 17490 21364 17500
rect 21644 17490 21700 17500
rect 21420 16772 21476 16782
rect 20524 16146 20580 16156
rect 20748 16770 21476 16772
rect 20748 16718 21422 16770
rect 21474 16718 21476 16770
rect 20748 16716 21476 16718
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19348 15372 19460 15428
rect 19740 15428 19796 15438
rect 19292 15362 19348 15372
rect 19740 15334 19796 15372
rect 20748 15426 20804 16716
rect 21420 16706 21476 16716
rect 21532 16772 21588 16782
rect 20748 15374 20750 15426
rect 20802 15374 20804 15426
rect 20748 15362 20804 15374
rect 20636 15090 20692 15102
rect 20636 15038 20638 15090
rect 20690 15038 20692 15090
rect 20636 14532 20692 15038
rect 20636 14466 20692 14476
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 19628 13858 19684 13870
rect 19628 13806 19630 13858
rect 19682 13806 19684 13858
rect 19516 13636 19572 13646
rect 19516 13542 19572 13580
rect 19404 13524 19460 13534
rect 19404 13430 19460 13468
rect 18844 11330 18900 11340
rect 19068 12348 19236 12404
rect 16604 11170 16996 11172
rect 16604 11118 16606 11170
rect 16658 11118 16996 11170
rect 16604 11116 16996 11118
rect 16604 11106 16660 11116
rect 15932 9998 15934 10050
rect 15986 9998 15988 10050
rect 15932 9986 15988 9998
rect 16044 9716 16100 9726
rect 16044 9714 16548 9716
rect 16044 9662 16046 9714
rect 16098 9662 16548 9714
rect 16044 9660 16548 9662
rect 16044 9650 16100 9660
rect 15484 9538 15540 9548
rect 14364 9102 14366 9154
rect 14418 9102 14420 9154
rect 14364 9090 14420 9102
rect 16492 8930 16548 9660
rect 16716 9604 16772 9614
rect 16716 9510 16772 9548
rect 16492 8878 16494 8930
rect 16546 8878 16548 8930
rect 16492 8866 16548 8878
rect 16828 8484 16884 8494
rect 16940 8484 16996 11116
rect 19068 10836 19124 12348
rect 19628 12292 19684 13806
rect 20300 13748 20356 13758
rect 20300 13654 20356 13692
rect 21532 13746 21588 16716
rect 21644 16660 21700 16670
rect 21644 16210 21700 16604
rect 21644 16158 21646 16210
rect 21698 16158 21700 16210
rect 21644 16146 21700 16158
rect 21756 14084 21812 17500
rect 22204 16660 22260 18956
rect 22316 18946 22372 18956
rect 22540 19012 22596 19022
rect 22540 18918 22596 18956
rect 22764 18338 22820 19070
rect 22876 19122 22932 19134
rect 22876 19070 22878 19122
rect 22930 19070 22932 19122
rect 22876 18564 22932 19070
rect 22876 18498 22932 18508
rect 22764 18286 22766 18338
rect 22818 18286 22820 18338
rect 22764 18274 22820 18286
rect 23212 18338 23268 19182
rect 23212 18286 23214 18338
rect 23266 18286 23268 18338
rect 22876 17668 22932 17678
rect 22316 16772 22372 16782
rect 22316 16678 22372 16716
rect 22204 16594 22260 16604
rect 22652 16660 22708 16670
rect 22652 16098 22708 16604
rect 22652 16046 22654 16098
rect 22706 16046 22708 16098
rect 22652 15202 22708 16046
rect 22652 15150 22654 15202
rect 22706 15150 22708 15202
rect 22652 15138 22708 15150
rect 21532 13694 21534 13746
rect 21586 13694 21588 13746
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19180 12236 19684 12292
rect 19180 11956 19236 12236
rect 20748 12180 20804 12190
rect 19292 12068 19348 12078
rect 19292 12066 19908 12068
rect 19292 12014 19294 12066
rect 19346 12014 19908 12066
rect 19292 12012 19908 12014
rect 19292 12002 19348 12012
rect 19180 11862 19236 11900
rect 19852 11506 19908 12012
rect 19852 11454 19854 11506
rect 19906 11454 19908 11506
rect 19852 11442 19908 11454
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19068 10770 19124 10780
rect 20748 10834 20804 12124
rect 20748 10782 20750 10834
rect 20802 10782 20804 10834
rect 20748 10770 20804 10782
rect 21420 11732 21476 11742
rect 20972 10722 21028 10734
rect 20972 10670 20974 10722
rect 21026 10670 21028 10722
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 17388 9042 17444 9054
rect 17388 8990 17390 9042
rect 17442 8990 17444 9042
rect 17388 8484 17444 8990
rect 16884 8428 17444 8484
rect 18172 8930 18228 8942
rect 20300 8932 20356 8942
rect 18172 8878 18174 8930
rect 18226 8878 18228 8930
rect 16828 8418 16884 8428
rect 17052 8370 17108 8428
rect 17052 8318 17054 8370
rect 17106 8318 17108 8370
rect 17052 8306 17108 8318
rect 18172 8372 18228 8878
rect 20076 8876 20300 8932
rect 18172 8306 18228 8316
rect 19404 8372 19460 8382
rect 19404 8278 19460 8316
rect 19628 8260 19684 8270
rect 19516 8034 19572 8046
rect 19516 7982 19518 8034
rect 19570 7982 19572 8034
rect 19516 7700 19572 7982
rect 19516 7634 19572 7644
rect 14140 7522 14196 7532
rect 18284 7588 18340 7598
rect 14028 7364 14084 7374
rect 14028 7362 14308 7364
rect 14028 7310 14030 7362
rect 14082 7310 14308 7362
rect 14028 7308 14308 7310
rect 14028 7298 14084 7308
rect 13580 6626 13636 6636
rect 12124 5966 12126 6018
rect 12178 5966 12180 6018
rect 12124 5954 12180 5966
rect 11340 5854 11342 5906
rect 11394 5854 11396 5906
rect 11340 5842 11396 5854
rect 14252 5794 14308 7308
rect 16156 6804 16212 6814
rect 14252 5742 14254 5794
rect 14306 5742 14308 5794
rect 14252 5730 14308 5742
rect 14700 6692 14756 6702
rect 14700 6130 14756 6636
rect 15036 6692 15092 6702
rect 15036 6598 15092 6636
rect 15372 6692 15428 6702
rect 15372 6598 15428 6636
rect 16156 6690 16212 6748
rect 18284 6802 18340 7532
rect 19628 7588 19684 8204
rect 20076 8258 20132 8876
rect 20300 8838 20356 8876
rect 20076 8206 20078 8258
rect 20130 8206 20132 8258
rect 20076 8194 20132 8206
rect 20188 8484 20244 8494
rect 19740 8148 19796 8158
rect 19740 8054 19796 8092
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 20076 7700 20132 7710
rect 20188 7700 20244 8428
rect 20972 8484 21028 10670
rect 21084 10610 21140 10622
rect 21084 10558 21086 10610
rect 21138 10558 21140 10610
rect 21084 9940 21140 10558
rect 21420 10050 21476 11676
rect 21532 11394 21588 13694
rect 21644 14028 21812 14084
rect 22876 14530 22932 17612
rect 23212 16660 23268 18286
rect 23548 17554 23604 19964
rect 23548 17502 23550 17554
rect 23602 17502 23604 17554
rect 23212 16594 23268 16604
rect 23324 17442 23380 17454
rect 23324 17390 23326 17442
rect 23378 17390 23380 17442
rect 23324 16324 23380 17390
rect 23548 16772 23604 17502
rect 23660 18564 23716 18574
rect 23660 17556 23716 18508
rect 23660 17462 23716 17500
rect 23548 16706 23604 16716
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 21644 11788 21700 14028
rect 22204 13634 22260 13646
rect 22204 13582 22206 13634
rect 22258 13582 22260 13634
rect 21868 13524 21924 13534
rect 21868 12964 21924 13468
rect 22204 13074 22260 13582
rect 22876 13524 22932 14478
rect 23212 16268 23380 16324
rect 22876 13458 22932 13468
rect 23100 14418 23156 14430
rect 23100 14366 23102 14418
rect 23154 14366 23156 14418
rect 22204 13022 22206 13074
rect 22258 13022 22260 13074
rect 22204 13010 22260 13022
rect 21756 12962 21924 12964
rect 21756 12910 21870 12962
rect 21922 12910 21924 12962
rect 21756 12908 21924 12910
rect 21756 12178 21812 12908
rect 21868 12898 21924 12908
rect 22092 12962 22148 12974
rect 22092 12910 22094 12962
rect 22146 12910 22148 12962
rect 22092 12292 22148 12910
rect 22428 12962 22484 12974
rect 22428 12910 22430 12962
rect 22482 12910 22484 12962
rect 22428 12852 22484 12910
rect 22428 12786 22484 12796
rect 22092 12236 22260 12292
rect 21756 12126 21758 12178
rect 21810 12126 21812 12178
rect 21756 12114 21812 12126
rect 21868 12180 21924 12190
rect 21868 12086 21924 12124
rect 22092 12066 22148 12078
rect 22092 12014 22094 12066
rect 22146 12014 22148 12066
rect 21644 11732 22036 11788
rect 21532 11342 21534 11394
rect 21586 11342 21588 11394
rect 21532 11172 21588 11342
rect 21532 11106 21588 11116
rect 21420 9998 21422 10050
rect 21474 9998 21476 10050
rect 21420 9986 21476 9998
rect 21980 10050 22036 11732
rect 22092 11508 22148 12014
rect 22204 11732 22260 12236
rect 22316 12180 22372 12190
rect 22316 12086 22372 12124
rect 22204 11666 22260 11676
rect 22204 11508 22260 11518
rect 22092 11506 22260 11508
rect 22092 11454 22206 11506
rect 22258 11454 22260 11506
rect 22092 11452 22260 11454
rect 22204 11442 22260 11452
rect 21980 9998 21982 10050
rect 22034 9998 22036 10050
rect 21980 9986 22036 9998
rect 21308 9940 21364 9950
rect 21084 9884 21308 9940
rect 21308 9826 21364 9884
rect 21308 9774 21310 9826
rect 21362 9774 21364 9826
rect 21308 9762 21364 9774
rect 22092 9940 22148 9950
rect 22092 9826 22148 9884
rect 22092 9774 22094 9826
rect 22146 9774 22148 9826
rect 22092 9762 22148 9774
rect 22764 9940 22820 9950
rect 22764 9826 22820 9884
rect 22764 9774 22766 9826
rect 22818 9774 22820 9826
rect 22764 9762 22820 9774
rect 23100 9826 23156 14366
rect 23212 14420 23268 16268
rect 23436 15986 23492 15998
rect 23436 15934 23438 15986
rect 23490 15934 23492 15986
rect 23436 15148 23492 15934
rect 23324 15092 23492 15148
rect 23772 15148 23828 26852
rect 24108 26852 24164 28028
rect 24220 28018 24276 28028
rect 23884 25508 23940 25518
rect 23884 25414 23940 25452
rect 24108 25396 24164 26796
rect 24220 27748 24276 27758
rect 24220 27074 24276 27692
rect 24220 27022 24222 27074
rect 24274 27022 24276 27074
rect 24220 25618 24276 27022
rect 24220 25566 24222 25618
rect 24274 25566 24276 25618
rect 24220 25554 24276 25566
rect 24332 26962 24388 26974
rect 24332 26910 24334 26962
rect 24386 26910 24388 26962
rect 24108 25330 24164 25340
rect 24332 22372 24388 26910
rect 24332 22306 24388 22316
rect 23996 22148 24052 22158
rect 24332 22148 24388 22158
rect 24052 22146 24388 22148
rect 24052 22094 24334 22146
rect 24386 22094 24388 22146
rect 24052 22092 24388 22094
rect 23996 22054 24052 22092
rect 24332 22082 24388 22092
rect 23884 21700 23940 21710
rect 23884 21606 23940 21644
rect 23996 19908 24052 19918
rect 23996 19346 24052 19852
rect 23996 19294 23998 19346
rect 24050 19294 24052 19346
rect 23996 19282 24052 19294
rect 24108 16882 24164 16894
rect 24108 16830 24110 16882
rect 24162 16830 24164 16882
rect 24108 15314 24164 16830
rect 24108 15262 24110 15314
rect 24162 15262 24164 15314
rect 23772 15092 23940 15148
rect 23324 14642 23380 15092
rect 23324 14590 23326 14642
rect 23378 14590 23380 14642
rect 23324 14578 23380 14590
rect 23436 14420 23492 14430
rect 23212 14418 23492 14420
rect 23212 14366 23438 14418
rect 23490 14366 23492 14418
rect 23212 14364 23492 14366
rect 23436 14354 23492 14364
rect 23884 12628 23940 15092
rect 24108 15092 24164 15262
rect 24444 15148 24500 31276
rect 24556 31276 24724 31332
rect 24556 31108 24612 31276
rect 24556 31042 24612 31052
rect 24668 30996 24724 31006
rect 24668 30902 24724 30940
rect 24556 29988 24612 29998
rect 24556 29894 24612 29932
rect 24668 27300 24724 27310
rect 24668 27186 24724 27244
rect 24668 27134 24670 27186
rect 24722 27134 24724 27186
rect 24668 27122 24724 27134
rect 24556 25508 24612 25518
rect 24556 25414 24612 25452
rect 24668 24948 24724 24958
rect 24668 24050 24724 24892
rect 24668 23998 24670 24050
rect 24722 23998 24724 24050
rect 24668 23986 24724 23998
rect 24668 22146 24724 22158
rect 24668 22094 24670 22146
rect 24722 22094 24724 22146
rect 24668 21924 24724 22094
rect 24668 21858 24724 21868
rect 24780 21588 24836 33964
rect 25228 31668 25284 37100
rect 25340 37090 25396 37100
rect 26908 36932 26964 36942
rect 26964 36876 27076 36932
rect 26908 36866 26964 36876
rect 25340 34914 25396 34926
rect 25340 34862 25342 34914
rect 25394 34862 25396 34914
rect 25340 32116 25396 34862
rect 26124 34804 26180 34814
rect 25788 34802 26180 34804
rect 25788 34750 26126 34802
rect 26178 34750 26180 34802
rect 25788 34748 26180 34750
rect 25452 34692 25508 34702
rect 25452 34130 25508 34636
rect 25788 34354 25844 34748
rect 26124 34738 26180 34748
rect 25788 34302 25790 34354
rect 25842 34302 25844 34354
rect 25788 34290 25844 34302
rect 25452 34078 25454 34130
rect 25506 34078 25508 34130
rect 25452 34066 25508 34078
rect 25900 34130 25956 34142
rect 25900 34078 25902 34130
rect 25954 34078 25956 34130
rect 25900 33346 25956 34078
rect 26012 34130 26068 34142
rect 26012 34078 26014 34130
rect 26066 34078 26068 34130
rect 26012 34020 26068 34078
rect 26012 33954 26068 33964
rect 25900 33294 25902 33346
rect 25954 33294 25956 33346
rect 25900 33282 25956 33294
rect 25564 33234 25620 33246
rect 25564 33182 25566 33234
rect 25618 33182 25620 33234
rect 25564 32900 25620 33182
rect 25676 33124 25732 33134
rect 26348 33124 26404 33134
rect 25676 33122 26404 33124
rect 25676 33070 25678 33122
rect 25730 33070 26350 33122
rect 26402 33070 26404 33122
rect 25676 33068 26404 33070
rect 25676 33058 25732 33068
rect 25564 32844 25844 32900
rect 25452 32788 25508 32798
rect 25508 32732 25732 32788
rect 25452 32722 25508 32732
rect 25676 32674 25732 32732
rect 25676 32622 25678 32674
rect 25730 32622 25732 32674
rect 25676 32610 25732 32622
rect 25564 32450 25620 32462
rect 25564 32398 25566 32450
rect 25618 32398 25620 32450
rect 25340 31780 25396 32060
rect 25452 32338 25508 32350
rect 25452 32286 25454 32338
rect 25506 32286 25508 32338
rect 25452 32004 25508 32286
rect 25452 31938 25508 31948
rect 25452 31780 25508 31790
rect 25340 31778 25508 31780
rect 25340 31726 25454 31778
rect 25506 31726 25508 31778
rect 25340 31724 25508 31726
rect 25452 31714 25508 31724
rect 25228 31612 25396 31668
rect 25116 31554 25172 31566
rect 25116 31502 25118 31554
rect 25170 31502 25172 31554
rect 25004 31332 25060 31342
rect 25116 31332 25172 31502
rect 25060 31276 25172 31332
rect 25004 31266 25060 31276
rect 25116 31108 25172 31118
rect 25116 30322 25172 31052
rect 25228 30996 25284 31006
rect 25228 30902 25284 30940
rect 25116 30270 25118 30322
rect 25170 30270 25172 30322
rect 25116 30258 25172 30270
rect 25340 29876 25396 31612
rect 25340 29810 25396 29820
rect 25452 31556 25508 31566
rect 25228 29652 25284 29662
rect 25116 28980 25172 28990
rect 24892 28644 24948 28654
rect 24892 28550 24948 28588
rect 25004 27076 25060 27086
rect 25004 26982 25060 27020
rect 25116 22482 25172 28924
rect 25228 28866 25284 29596
rect 25228 28814 25230 28866
rect 25282 28814 25284 28866
rect 25228 28802 25284 28814
rect 25340 28644 25396 28654
rect 25340 28082 25396 28588
rect 25340 28030 25342 28082
rect 25394 28030 25396 28082
rect 25340 27074 25396 28030
rect 25340 27022 25342 27074
rect 25394 27022 25396 27074
rect 25228 26964 25284 27002
rect 25228 26898 25284 26908
rect 25340 26852 25396 27022
rect 25340 26786 25396 26796
rect 25452 27972 25508 31500
rect 25564 30994 25620 32398
rect 25788 31668 25844 32844
rect 26236 32788 26292 32798
rect 26236 32004 26292 32732
rect 26236 31938 26292 31948
rect 25788 31556 25844 31612
rect 26236 31666 26292 31678
rect 26236 31614 26238 31666
rect 26290 31614 26292 31666
rect 25788 31500 26068 31556
rect 26012 31106 26068 31500
rect 26012 31054 26014 31106
rect 26066 31054 26068 31106
rect 26012 31042 26068 31054
rect 25564 30942 25566 30994
rect 25618 30942 25620 30994
rect 25564 30930 25620 30942
rect 25788 30994 25844 31006
rect 25788 30942 25790 30994
rect 25842 30942 25844 30994
rect 25788 30884 25844 30942
rect 25788 30818 25844 30828
rect 25900 30884 25956 30894
rect 26236 30884 26292 31614
rect 25900 30882 26292 30884
rect 25900 30830 25902 30882
rect 25954 30830 26292 30882
rect 25900 30828 26292 30830
rect 25900 30818 25956 30828
rect 25564 30212 25620 30222
rect 25564 28866 25620 30156
rect 26236 30212 26292 30222
rect 26236 30118 26292 30156
rect 26124 29316 26180 29326
rect 26124 29222 26180 29260
rect 25564 28814 25566 28866
rect 25618 28814 25620 28866
rect 25564 28644 25620 28814
rect 25788 28756 25844 28766
rect 25788 28662 25844 28700
rect 26236 28756 26292 28766
rect 25564 28578 25620 28588
rect 26236 28642 26292 28700
rect 26236 28590 26238 28642
rect 26290 28590 26292 28642
rect 26236 28578 26292 28590
rect 25228 25396 25284 25406
rect 25228 25302 25284 25340
rect 25228 23716 25284 23726
rect 25228 23622 25284 23660
rect 25116 22430 25118 22482
rect 25170 22430 25172 22482
rect 25116 22418 25172 22430
rect 24780 20132 24836 21532
rect 24780 20038 24836 20076
rect 25228 20018 25284 20030
rect 25228 19966 25230 20018
rect 25282 19966 25284 20018
rect 25228 18900 25284 19966
rect 25340 19908 25396 19918
rect 25340 19814 25396 19852
rect 25116 18844 25284 18900
rect 25116 18674 25172 18844
rect 25452 18788 25508 27916
rect 25676 28420 25732 28430
rect 25676 27076 25732 28364
rect 26236 27746 26292 27758
rect 26236 27694 26238 27746
rect 26290 27694 26292 27746
rect 25676 26516 25732 27020
rect 25788 27076 25844 27086
rect 26236 27076 26292 27694
rect 25788 27074 26292 27076
rect 25788 27022 25790 27074
rect 25842 27022 26292 27074
rect 25788 27020 26292 27022
rect 25788 26852 25844 27020
rect 25788 26786 25844 26796
rect 25788 26516 25844 26526
rect 25676 26514 25844 26516
rect 25676 26462 25790 26514
rect 25842 26462 25844 26514
rect 25676 26460 25844 26462
rect 25788 26450 25844 26460
rect 26236 26516 26292 27020
rect 26236 26450 26292 26460
rect 26348 25844 26404 33068
rect 26460 30884 26516 30894
rect 26516 30828 26628 30884
rect 26460 30790 26516 30828
rect 26460 29316 26516 29326
rect 26460 28980 26516 29260
rect 26460 28914 26516 28924
rect 26460 28644 26516 28654
rect 26460 28418 26516 28588
rect 26460 28366 26462 28418
rect 26514 28366 26516 28418
rect 26460 26964 26516 28366
rect 26460 26898 26516 26908
rect 26124 25788 26404 25844
rect 25564 25506 25620 25518
rect 25564 25454 25566 25506
rect 25618 25454 25620 25506
rect 25564 24948 25620 25454
rect 25564 24882 25620 24892
rect 25788 25508 25844 25518
rect 25788 24948 25844 25452
rect 25788 24854 25844 24892
rect 26012 25394 26068 25406
rect 26012 25342 26014 25394
rect 26066 25342 26068 25394
rect 25676 23938 25732 23950
rect 25676 23886 25678 23938
rect 25730 23886 25732 23938
rect 25676 23492 25732 23886
rect 25676 23426 25732 23436
rect 25564 22146 25620 22158
rect 25564 22094 25566 22146
rect 25618 22094 25620 22146
rect 25564 21924 25620 22094
rect 25900 22148 25956 22158
rect 25900 22054 25956 22092
rect 25564 21858 25620 21868
rect 25788 20132 25844 20142
rect 25788 20038 25844 20076
rect 25564 20020 25620 20030
rect 25564 19926 25620 19964
rect 25116 18622 25118 18674
rect 25170 18622 25172 18674
rect 25116 18610 25172 18622
rect 25228 18732 25508 18788
rect 26012 19348 26068 25342
rect 26124 24052 26180 25788
rect 26348 25620 26404 25630
rect 26348 25526 26404 25564
rect 26236 25506 26292 25518
rect 26236 25454 26238 25506
rect 26290 25454 26292 25506
rect 26236 24724 26292 25454
rect 26236 24610 26292 24668
rect 26236 24558 26238 24610
rect 26290 24558 26292 24610
rect 26236 24546 26292 24558
rect 26124 23958 26180 23996
rect 26124 23716 26180 23726
rect 26124 23044 26180 23660
rect 26460 23154 26516 23166
rect 26460 23102 26462 23154
rect 26514 23102 26516 23154
rect 26460 23044 26516 23102
rect 26124 23042 26516 23044
rect 26124 22990 26126 23042
rect 26178 22990 26516 23042
rect 26124 22988 26516 22990
rect 26124 22978 26180 22988
rect 26124 19348 26180 19358
rect 26012 19346 26180 19348
rect 26012 19294 26126 19346
rect 26178 19294 26180 19346
rect 26012 19292 26180 19294
rect 25228 17220 25284 18732
rect 25340 18564 25396 18574
rect 25340 18470 25396 18508
rect 26012 18564 26068 19292
rect 26124 19282 26180 19292
rect 26012 18498 26068 18508
rect 25116 17164 25284 17220
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 25452 17556 25508 18398
rect 26236 18450 26292 22988
rect 26460 22484 26516 22494
rect 26572 22484 26628 30828
rect 26908 28756 26964 28766
rect 26908 28662 26964 28700
rect 26908 28084 26964 28094
rect 27020 28084 27076 36876
rect 27132 34244 27188 37100
rect 27132 34178 27188 34188
rect 27356 29876 27412 29886
rect 27356 28756 27412 29820
rect 27356 28662 27412 28700
rect 26908 28082 27300 28084
rect 26908 28030 26910 28082
rect 26962 28030 27300 28082
rect 26908 28028 27300 28030
rect 26908 28018 26964 28028
rect 27244 27858 27300 28028
rect 27244 27806 27246 27858
rect 27298 27806 27300 27858
rect 27244 27794 27300 27806
rect 27468 27636 27524 38612
rect 28140 38050 28196 43260
rect 28588 43250 28644 43260
rect 29036 43314 29092 43326
rect 29036 43262 29038 43314
rect 29090 43262 29092 43314
rect 28588 42532 28644 42542
rect 29036 42532 29092 43262
rect 28588 42530 29092 42532
rect 28588 42478 28590 42530
rect 28642 42478 29092 42530
rect 28588 42476 29092 42478
rect 28588 40740 28644 42476
rect 28588 40674 28644 40684
rect 29148 41970 29204 44270
rect 30156 45444 30212 45454
rect 29932 44212 29988 44222
rect 29372 44210 29988 44212
rect 29372 44158 29934 44210
rect 29986 44158 29988 44210
rect 29372 44156 29988 44158
rect 29372 43762 29428 44156
rect 29932 44146 29988 44156
rect 29372 43710 29374 43762
rect 29426 43710 29428 43762
rect 29372 43698 29428 43710
rect 29260 43540 29316 43550
rect 29260 43446 29316 43484
rect 29708 43428 29764 43438
rect 29372 43316 29428 43326
rect 29372 43222 29428 43260
rect 29708 42978 29764 43372
rect 29708 42926 29710 42978
rect 29762 42926 29764 42978
rect 29708 42914 29764 42926
rect 29820 42530 29876 42542
rect 29820 42478 29822 42530
rect 29874 42478 29876 42530
rect 29820 42082 29876 42478
rect 29932 42530 29988 42542
rect 29932 42478 29934 42530
rect 29986 42478 29988 42530
rect 29932 42420 29988 42478
rect 30044 42420 30100 42430
rect 29932 42364 30044 42420
rect 30044 42354 30100 42364
rect 29820 42030 29822 42082
rect 29874 42030 29876 42082
rect 29820 42018 29876 42030
rect 29148 41918 29150 41970
rect 29202 41918 29204 41970
rect 29148 41300 29204 41918
rect 29148 40404 29204 41244
rect 29148 40310 29204 40348
rect 28700 40290 28756 40302
rect 28700 40238 28702 40290
rect 28754 40238 28756 40290
rect 28364 39620 28420 39630
rect 28700 39620 28756 40238
rect 28364 39618 28756 39620
rect 28364 39566 28366 39618
rect 28418 39566 28756 39618
rect 28364 39564 28756 39566
rect 28364 38668 28420 39564
rect 30044 38836 30100 38846
rect 30156 38836 30212 45388
rect 30044 38834 30212 38836
rect 30044 38782 30046 38834
rect 30098 38782 30212 38834
rect 30044 38780 30212 38782
rect 30044 38770 30100 38780
rect 29260 38724 29316 38762
rect 29596 38724 29652 38734
rect 29260 38722 29652 38724
rect 29260 38670 29262 38722
rect 29314 38670 29598 38722
rect 29650 38670 29652 38722
rect 29260 38668 29652 38670
rect 28140 37998 28142 38050
rect 28194 37998 28196 38050
rect 28140 37986 28196 37998
rect 28252 38612 28420 38668
rect 29036 38612 29316 38668
rect 29596 38658 29652 38668
rect 30268 38668 30324 46396
rect 30940 45444 30996 46734
rect 30940 45378 30996 45388
rect 32284 45332 32340 45342
rect 32060 45106 32116 45118
rect 32060 45054 32062 45106
rect 32114 45054 32116 45106
rect 31500 44996 31556 45006
rect 31500 44902 31556 44940
rect 32060 44436 32116 45054
rect 32284 45106 32340 45276
rect 32284 45054 32286 45106
rect 32338 45054 32340 45106
rect 32284 45042 32340 45054
rect 32060 44342 32116 44380
rect 32508 44434 32564 46844
rect 33516 46788 33572 46798
rect 33516 46694 33572 46732
rect 33740 46676 33796 47516
rect 35308 47572 35364 47582
rect 35308 47478 35364 47516
rect 33628 46674 33796 46676
rect 33628 46622 33742 46674
rect 33794 46622 33796 46674
rect 33628 46620 33796 46622
rect 33628 45444 33684 46620
rect 33740 46610 33796 46620
rect 35532 47236 35588 48748
rect 36876 48804 36932 48814
rect 37100 48804 37156 50318
rect 37772 50036 37828 50046
rect 37772 50034 38276 50036
rect 37772 49982 37774 50034
rect 37826 49982 38276 50034
rect 37772 49980 38276 49982
rect 37772 49970 37828 49980
rect 37436 49812 37492 49822
rect 37436 49718 37492 49756
rect 37548 49810 37604 49822
rect 37548 49758 37550 49810
rect 37602 49758 37604 49810
rect 36932 48802 37156 48804
rect 36932 48750 37102 48802
rect 37154 48750 37156 48802
rect 36932 48748 37156 48750
rect 36876 48738 36932 48748
rect 37100 47572 37156 48748
rect 37100 47506 37156 47516
rect 37212 48916 37268 48926
rect 35756 47236 35812 47246
rect 35532 47234 35812 47236
rect 35532 47182 35758 47234
rect 35810 47182 35812 47234
rect 35532 47180 35812 47182
rect 35532 46674 35588 47180
rect 35756 47170 35812 47180
rect 35532 46622 35534 46674
rect 35586 46622 35588 46674
rect 35532 46610 35588 46622
rect 36204 46564 36260 46574
rect 36204 46470 36260 46508
rect 37100 46564 37156 46574
rect 35196 46284 35460 46294
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35196 46218 35460 46228
rect 37100 46002 37156 46508
rect 37100 45950 37102 46002
rect 37154 45950 37156 46002
rect 37100 45938 37156 45950
rect 33964 45892 34020 45902
rect 33964 45890 34244 45892
rect 33964 45838 33966 45890
rect 34018 45838 34244 45890
rect 33964 45836 34244 45838
rect 33964 45826 34020 45836
rect 33516 45388 33684 45444
rect 34076 45666 34132 45678
rect 34076 45614 34078 45666
rect 34130 45614 34132 45666
rect 33404 45218 33460 45230
rect 33404 45166 33406 45218
rect 33458 45166 33460 45218
rect 32508 44382 32510 44434
rect 32562 44382 32564 44434
rect 32508 44370 32564 44382
rect 32844 44996 32900 45006
rect 32844 44436 32900 44940
rect 33292 44884 33348 44894
rect 33292 44790 33348 44828
rect 32844 44342 32900 44380
rect 33404 44436 33460 45166
rect 33516 44996 33572 45388
rect 34076 45332 34132 45614
rect 33628 45276 34132 45332
rect 33628 45218 33684 45276
rect 33628 45166 33630 45218
rect 33682 45166 33684 45218
rect 33628 45154 33684 45166
rect 33516 44940 33684 44996
rect 33404 44370 33460 44380
rect 32956 44100 33012 44110
rect 33404 44100 33460 44110
rect 32956 44098 33460 44100
rect 32956 44046 32958 44098
rect 33010 44046 33406 44098
rect 33458 44046 33460 44098
rect 32956 44044 33460 44046
rect 32956 42756 33012 44044
rect 33404 44034 33460 44044
rect 33516 43538 33572 43550
rect 33516 43486 33518 43538
rect 33570 43486 33572 43538
rect 33068 42756 33124 42766
rect 32956 42754 33124 42756
rect 32956 42702 33070 42754
rect 33122 42702 33124 42754
rect 32956 42700 33124 42702
rect 30492 42530 30548 42542
rect 32284 42532 32340 42542
rect 32732 42532 32788 42542
rect 30492 42478 30494 42530
rect 30546 42478 30548 42530
rect 30492 42420 30548 42478
rect 30492 42354 30548 42364
rect 32172 42530 32732 42532
rect 32172 42478 32286 42530
rect 32338 42478 32732 42530
rect 32172 42476 32732 42478
rect 31948 41860 32004 41870
rect 31948 40402 32004 41804
rect 32172 41636 32228 42476
rect 32284 42466 32340 42476
rect 32732 42438 32788 42476
rect 33068 41972 33124 42700
rect 33292 42754 33348 42766
rect 33292 42702 33294 42754
rect 33346 42702 33348 42754
rect 33292 42532 33348 42702
rect 33292 42466 33348 42476
rect 33516 42754 33572 43486
rect 33628 43540 33684 44940
rect 34188 44994 34244 45836
rect 34300 45890 34356 45902
rect 34300 45838 34302 45890
rect 34354 45838 34356 45890
rect 34300 45108 34356 45838
rect 36988 45780 37044 45790
rect 36876 45724 36988 45780
rect 36316 45668 36372 45678
rect 34860 45220 34916 45230
rect 34636 45108 34692 45118
rect 34300 45052 34636 45108
rect 34692 45052 34804 45108
rect 34636 45014 34692 45052
rect 34188 44942 34190 44994
rect 34242 44942 34244 44994
rect 33964 44436 34020 44446
rect 33964 44342 34020 44380
rect 34188 44324 34244 44942
rect 34300 44884 34356 44894
rect 34300 44790 34356 44828
rect 34748 44324 34804 45052
rect 33740 43764 33796 43774
rect 33740 43670 33796 43708
rect 34188 43764 34244 44268
rect 34188 43698 34244 43708
rect 34412 44322 34804 44324
rect 34412 44270 34750 44322
rect 34802 44270 34804 44322
rect 34412 44268 34804 44270
rect 34412 43762 34468 44268
rect 34748 44258 34804 44268
rect 34860 44436 34916 45164
rect 35420 45108 35476 45118
rect 35644 45108 35700 45118
rect 35420 45106 35700 45108
rect 35420 45054 35422 45106
rect 35474 45054 35646 45106
rect 35698 45054 35700 45106
rect 35420 45052 35700 45054
rect 35420 44996 35476 45052
rect 35644 45042 35700 45052
rect 35756 45108 35812 45118
rect 35756 45014 35812 45052
rect 35420 44930 35476 44940
rect 36204 44882 36260 44894
rect 36204 44830 36206 44882
rect 36258 44830 36260 44882
rect 35196 44716 35460 44726
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35196 44650 35460 44660
rect 34860 44210 34916 44380
rect 35756 44324 35812 44334
rect 36204 44324 36260 44830
rect 35812 44268 36260 44324
rect 35756 44230 35812 44268
rect 34860 44158 34862 44210
rect 34914 44158 34916 44210
rect 34860 44146 34916 44158
rect 36316 44098 36372 45612
rect 36540 45332 36596 45342
rect 36876 45332 36932 45724
rect 36988 45686 37044 45724
rect 37212 45556 37268 48860
rect 37548 48916 37604 49758
rect 37884 49810 37940 49822
rect 37884 49758 37886 49810
rect 37938 49758 37940 49810
rect 37660 49698 37716 49710
rect 37660 49646 37662 49698
rect 37714 49646 37716 49698
rect 37660 49476 37716 49646
rect 37660 49410 37716 49420
rect 37884 49476 37940 49758
rect 37884 49028 37940 49420
rect 37548 48850 37604 48860
rect 37660 48972 37940 49028
rect 38220 49028 38276 49980
rect 38444 50034 38500 50428
rect 38444 49982 38446 50034
rect 38498 49982 38500 50034
rect 38444 49970 38500 49982
rect 38556 49812 38612 49822
rect 38332 49586 38388 49598
rect 38332 49534 38334 49586
rect 38386 49534 38388 49586
rect 38332 49138 38388 49534
rect 38332 49086 38334 49138
rect 38386 49086 38388 49138
rect 38332 49074 38388 49086
rect 37548 46452 37604 46462
rect 37548 45890 37604 46396
rect 37548 45838 37550 45890
rect 37602 45838 37604 45890
rect 37548 45826 37604 45838
rect 36540 45330 36932 45332
rect 36540 45278 36542 45330
rect 36594 45278 36932 45330
rect 36540 45276 36932 45278
rect 36988 45500 37268 45556
rect 37324 45778 37380 45790
rect 37324 45726 37326 45778
rect 37378 45726 37380 45778
rect 36540 45266 36596 45276
rect 36316 44046 36318 44098
rect 36370 44046 36372 44098
rect 36316 44034 36372 44046
rect 36428 44882 36484 44894
rect 36428 44830 36430 44882
rect 36482 44830 36484 44882
rect 36428 44210 36484 44830
rect 36988 44884 37044 45500
rect 37324 45332 37380 45726
rect 37324 45238 37380 45276
rect 37100 45108 37156 45118
rect 37436 45108 37492 45118
rect 37100 45106 37436 45108
rect 37100 45054 37102 45106
rect 37154 45054 37436 45106
rect 37100 45052 37436 45054
rect 37100 45042 37156 45052
rect 37436 45014 37492 45052
rect 36988 44828 37156 44884
rect 36428 44158 36430 44210
rect 36482 44158 36484 44210
rect 34412 43710 34414 43762
rect 34466 43710 34468 43762
rect 34412 43698 34468 43710
rect 33964 43540 34020 43550
rect 33628 43484 33796 43540
rect 33516 42702 33518 42754
rect 33570 42702 33572 42754
rect 33180 42196 33236 42206
rect 33516 42196 33572 42702
rect 33516 42140 33684 42196
rect 33180 42102 33236 42140
rect 33516 41972 33572 41982
rect 33068 41970 33572 41972
rect 33068 41918 33518 41970
rect 33570 41918 33572 41970
rect 33068 41916 33572 41918
rect 33516 41906 33572 41916
rect 33180 41746 33236 41758
rect 33180 41694 33182 41746
rect 33234 41694 33236 41746
rect 33180 41636 33236 41694
rect 33292 41748 33348 41758
rect 33628 41748 33684 42140
rect 33292 41654 33348 41692
rect 33404 41692 33684 41748
rect 32172 41570 32228 41580
rect 32284 41580 33236 41636
rect 31948 40350 31950 40402
rect 32002 40350 32004 40402
rect 31948 40338 32004 40350
rect 32172 40402 32228 40414
rect 32172 40350 32174 40402
rect 32226 40350 32228 40402
rect 32172 40292 32228 40350
rect 32172 40226 32228 40236
rect 30940 38946 30996 38958
rect 30940 38894 30942 38946
rect 30994 38894 30996 38946
rect 30492 38836 30548 38846
rect 30828 38836 30884 38846
rect 30492 38834 30884 38836
rect 30492 38782 30494 38834
rect 30546 38782 30830 38834
rect 30882 38782 30884 38834
rect 30492 38780 30884 38782
rect 30492 38770 30548 38780
rect 30828 38770 30884 38780
rect 30940 38668 30996 38894
rect 32060 38722 32116 38734
rect 32060 38670 32062 38722
rect 32114 38670 32116 38722
rect 30268 38612 30772 38668
rect 30940 38612 31444 38668
rect 28028 37380 28084 37390
rect 28028 37286 28084 37324
rect 28140 36484 28196 36494
rect 28252 36484 28308 38612
rect 28476 38050 28532 38062
rect 28476 37998 28478 38050
rect 28530 37998 28532 38050
rect 28476 37828 28532 37998
rect 28588 37940 28644 37950
rect 28588 37846 28644 37884
rect 28476 37492 28532 37772
rect 28476 37436 28868 37492
rect 28476 37266 28532 37278
rect 28476 37214 28478 37266
rect 28530 37214 28532 37266
rect 28476 36596 28532 37214
rect 28588 36596 28644 36606
rect 28476 36594 28644 36596
rect 28476 36542 28590 36594
rect 28642 36542 28644 36594
rect 28476 36540 28644 36542
rect 28588 36530 28644 36540
rect 28140 36482 28308 36484
rect 28140 36430 28142 36482
rect 28194 36430 28308 36482
rect 28140 36428 28308 36430
rect 28364 36482 28420 36494
rect 28364 36430 28366 36482
rect 28418 36430 28420 36482
rect 28140 36418 28196 36428
rect 28364 36260 28420 36430
rect 28476 36260 28532 36270
rect 28364 36204 28476 36260
rect 28476 36194 28532 36204
rect 28140 36148 28196 36158
rect 28140 28868 28196 36092
rect 28700 35252 28756 35262
rect 28364 35026 28420 35038
rect 28364 34974 28366 35026
rect 28418 34974 28420 35026
rect 28364 34916 28420 34974
rect 28364 34850 28420 34860
rect 28700 34354 28756 35196
rect 28700 34302 28702 34354
rect 28754 34302 28756 34354
rect 28700 34290 28756 34302
rect 28364 32004 28420 32014
rect 28364 31890 28420 31948
rect 28364 31838 28366 31890
rect 28418 31838 28420 31890
rect 28364 31780 28420 31838
rect 28364 31714 28420 31724
rect 28140 28802 28196 28812
rect 28252 31668 28308 31678
rect 28252 28084 28308 31612
rect 28364 29314 28420 29326
rect 28364 29262 28366 29314
rect 28418 29262 28420 29314
rect 28364 28868 28420 29262
rect 28812 29204 28868 37436
rect 28924 37268 28980 37278
rect 28924 37174 28980 37212
rect 28924 29204 28980 29214
rect 28812 29148 28924 29204
rect 28364 28802 28420 28812
rect 28700 28532 28756 28542
rect 28252 28018 28308 28028
rect 28588 28476 28700 28532
rect 27468 27188 27524 27580
rect 27468 27122 27524 27132
rect 28588 27524 28644 28476
rect 28700 28466 28756 28476
rect 28588 26964 28644 27468
rect 28588 26898 28644 26908
rect 28700 27412 28756 27422
rect 28028 26180 28084 26190
rect 28028 26086 28084 26124
rect 28700 25172 28756 27356
rect 28812 26628 28868 26638
rect 28812 26290 28868 26572
rect 28924 26404 28980 29148
rect 29036 28532 29092 38612
rect 30044 38052 30100 38062
rect 30492 38052 30548 38062
rect 30044 38050 30548 38052
rect 30044 37998 30046 38050
rect 30098 37998 30494 38050
rect 30546 37998 30548 38050
rect 30044 37996 30548 37998
rect 30044 37986 30100 37996
rect 29484 37940 29540 37950
rect 29260 37828 29316 37838
rect 29260 37734 29316 37772
rect 29372 37492 29428 37502
rect 29372 37398 29428 37436
rect 29484 37378 29540 37884
rect 29484 37326 29486 37378
rect 29538 37326 29540 37378
rect 29484 37314 29540 37326
rect 30268 36482 30324 36494
rect 30268 36430 30270 36482
rect 30322 36430 30324 36482
rect 29148 36260 29204 36270
rect 29260 36260 29316 36270
rect 29204 36258 29316 36260
rect 29204 36206 29262 36258
rect 29314 36206 29316 36258
rect 29204 36204 29316 36206
rect 29148 35028 29204 36204
rect 29260 36194 29316 36204
rect 30268 35364 30324 36430
rect 30268 35298 30324 35308
rect 29148 33124 29204 34972
rect 29148 33058 29204 33068
rect 29260 35252 29316 35262
rect 29260 34914 29316 35196
rect 29260 34862 29262 34914
rect 29314 34862 29316 34914
rect 29260 32116 29316 34862
rect 29932 34804 29988 34814
rect 29932 34802 30212 34804
rect 29932 34750 29934 34802
rect 29986 34750 30212 34802
rect 29932 34748 30212 34750
rect 29932 34738 29988 34748
rect 29596 33572 29652 33582
rect 29596 33570 29876 33572
rect 29596 33518 29598 33570
rect 29650 33518 29876 33570
rect 29596 33516 29876 33518
rect 29596 33506 29652 33516
rect 29708 33348 29764 33358
rect 29820 33348 29876 33516
rect 30156 33570 30212 34748
rect 30380 34244 30436 34254
rect 30156 33518 30158 33570
rect 30210 33518 30212 33570
rect 30156 33506 30212 33518
rect 30268 34130 30324 34142
rect 30268 34078 30270 34130
rect 30322 34078 30324 34130
rect 29932 33348 29988 33358
rect 29820 33346 29988 33348
rect 29820 33294 29934 33346
rect 29986 33294 29988 33346
rect 29820 33292 29988 33294
rect 29708 33254 29764 33292
rect 29932 33282 29988 33292
rect 30268 33348 30324 34078
rect 30380 33908 30436 34188
rect 30380 33842 30436 33852
rect 30492 33348 30548 37996
rect 30716 38050 30772 38612
rect 31388 38162 31444 38612
rect 31388 38110 31390 38162
rect 31442 38110 31444 38162
rect 31388 38098 31444 38110
rect 30716 37998 30718 38050
rect 30770 37998 30772 38050
rect 30716 37986 30772 37998
rect 31948 37938 32004 37950
rect 31948 37886 31950 37938
rect 32002 37886 32004 37938
rect 31948 37492 32004 37886
rect 32060 37938 32116 38670
rect 32284 38050 32340 41580
rect 33180 41524 33236 41580
rect 33404 41524 33460 41692
rect 33180 41468 33460 41524
rect 32396 41300 32452 41310
rect 32396 41206 32452 41244
rect 33516 41300 33572 41310
rect 33516 41186 33572 41244
rect 33516 41134 33518 41186
rect 33570 41134 33572 41186
rect 33516 41122 33572 41134
rect 33292 40402 33348 40414
rect 33292 40350 33294 40402
rect 33346 40350 33348 40402
rect 32396 40290 32452 40302
rect 32396 40238 32398 40290
rect 32450 40238 32452 40290
rect 32396 38946 32452 40238
rect 33292 40292 33348 40350
rect 33292 40226 33348 40236
rect 32396 38894 32398 38946
rect 32450 38894 32452 38946
rect 32396 38882 32452 38894
rect 32508 38836 32564 38846
rect 33292 38836 33348 38846
rect 32508 38834 33348 38836
rect 32508 38782 32510 38834
rect 32562 38782 33294 38834
rect 33346 38782 33348 38834
rect 32508 38780 33348 38782
rect 32508 38770 32564 38780
rect 33292 38770 33348 38780
rect 33740 38834 33796 43484
rect 33964 42978 34020 43484
rect 33964 42926 33966 42978
rect 34018 42926 34020 42978
rect 33964 42914 34020 42926
rect 34076 43538 34132 43550
rect 34076 43486 34078 43538
rect 34130 43486 34132 43538
rect 34076 43428 34132 43486
rect 34076 42532 34132 43372
rect 34860 43428 34916 43438
rect 34860 43334 34916 43372
rect 35196 43148 35460 43158
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35196 43082 35460 43092
rect 36428 42980 36484 44158
rect 36428 42914 36484 42924
rect 36988 43316 37044 43326
rect 36988 42756 37044 43260
rect 36988 42662 37044 42700
rect 37100 42642 37156 44828
rect 37100 42590 37102 42642
rect 37154 42590 37156 42642
rect 37100 42578 37156 42590
rect 37660 42642 37716 48972
rect 38220 48934 38276 48972
rect 38556 49028 38612 49756
rect 38668 49810 38724 49822
rect 38668 49758 38670 49810
rect 38722 49758 38724 49810
rect 38668 49140 38724 49758
rect 38668 49074 38724 49084
rect 39788 49140 39844 49150
rect 38556 48934 38612 48972
rect 37996 48916 38052 48926
rect 37996 48822 38052 48860
rect 38668 48916 38724 48926
rect 38444 48804 38500 48814
rect 38444 48710 38500 48748
rect 37996 48244 38052 48254
rect 37996 46116 38052 48188
rect 38556 47572 38612 47582
rect 38556 47478 38612 47516
rect 38668 46898 38724 48860
rect 38668 46846 38670 46898
rect 38722 46846 38724 46898
rect 38332 46564 38388 46574
rect 38332 46470 38388 46508
rect 37996 46060 38612 46116
rect 37884 45780 37940 45790
rect 37884 45686 37940 45724
rect 37996 45778 38052 46060
rect 38556 46002 38612 46060
rect 38556 45950 38558 46002
rect 38610 45950 38612 46002
rect 38556 45938 38612 45950
rect 38220 45892 38276 45902
rect 38220 45798 38276 45836
rect 37996 45726 37998 45778
rect 38050 45726 38052 45778
rect 37996 45330 38052 45726
rect 38668 45780 38724 46846
rect 39004 48804 39060 48814
rect 38892 46676 38948 46686
rect 38892 46582 38948 46620
rect 38780 46564 38836 46574
rect 38780 46470 38836 46508
rect 38668 45714 38724 45724
rect 37996 45278 37998 45330
rect 38050 45278 38052 45330
rect 37996 45266 38052 45278
rect 38780 45332 38836 45342
rect 38332 45220 38388 45230
rect 38332 45126 38388 45164
rect 38444 45108 38500 45118
rect 38444 44100 38500 45052
rect 38780 45106 38836 45276
rect 38892 45220 38948 45230
rect 38892 45126 38948 45164
rect 38780 45054 38782 45106
rect 38834 45054 38836 45106
rect 38780 45042 38836 45054
rect 38668 44100 38724 44110
rect 38444 44044 38668 44100
rect 38668 44006 38724 44044
rect 38892 43764 38948 43774
rect 39004 43764 39060 48748
rect 39788 48466 39844 49084
rect 39788 48414 39790 48466
rect 39842 48414 39844 48466
rect 39788 48402 39844 48414
rect 40012 49028 40068 49038
rect 40012 47460 40068 48972
rect 40348 48804 40404 50654
rect 40348 48738 40404 48748
rect 40124 48242 40180 48254
rect 40124 48190 40126 48242
rect 40178 48190 40180 48242
rect 40124 48132 40180 48190
rect 40124 48066 40180 48076
rect 40012 46898 40068 47404
rect 40012 46846 40014 46898
rect 40066 46846 40068 46898
rect 40012 46834 40068 46846
rect 39340 46674 39396 46686
rect 39340 46622 39342 46674
rect 39394 46622 39396 46674
rect 39340 46564 39396 46622
rect 40012 46676 40068 46686
rect 39676 46564 39732 46574
rect 39340 46562 39732 46564
rect 39340 46510 39678 46562
rect 39730 46510 39732 46562
rect 39340 46508 39732 46510
rect 39564 45780 39620 45790
rect 39564 45686 39620 45724
rect 39452 45220 39508 45230
rect 39452 45126 39508 45164
rect 38892 43762 39060 43764
rect 38892 43710 38894 43762
rect 38946 43710 39060 43762
rect 38892 43708 39060 43710
rect 39564 44100 39620 44110
rect 38892 43698 38948 43708
rect 38780 43538 38836 43550
rect 38780 43486 38782 43538
rect 38834 43486 38836 43538
rect 38332 42980 38388 42990
rect 37772 42756 37828 42766
rect 37772 42662 37828 42700
rect 37660 42590 37662 42642
rect 37714 42590 37716 42642
rect 37660 42578 37716 42590
rect 34076 42466 34132 42476
rect 37324 42530 37380 42542
rect 37324 42478 37326 42530
rect 37378 42478 37380 42530
rect 36652 41858 36708 41870
rect 36652 41806 36654 41858
rect 36706 41806 36708 41858
rect 35196 41580 35460 41590
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35196 41514 35460 41524
rect 35756 41300 35812 41310
rect 34300 41076 34356 41086
rect 34300 40982 34356 41020
rect 35308 40516 35364 40526
rect 33740 38782 33742 38834
rect 33794 38782 33796 38834
rect 33740 38770 33796 38782
rect 34860 40460 35308 40516
rect 34860 39058 34916 40460
rect 35308 40422 35364 40460
rect 35756 40290 35812 41244
rect 35756 40238 35758 40290
rect 35810 40238 35812 40290
rect 35756 40226 35812 40238
rect 36428 41298 36484 41310
rect 36428 41246 36430 41298
rect 36482 41246 36484 41298
rect 35196 40012 35460 40022
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35196 39946 35460 39956
rect 36428 39620 36484 41246
rect 36652 41300 36708 41806
rect 36652 41234 36708 41244
rect 37324 41186 37380 42478
rect 37324 41134 37326 41186
rect 37378 41134 37380 41186
rect 37324 41122 37380 41134
rect 37436 42530 37492 42542
rect 37436 42478 37438 42530
rect 37490 42478 37492 42530
rect 36988 41074 37044 41086
rect 36988 41022 36990 41074
rect 37042 41022 37044 41074
rect 36988 39844 37044 41022
rect 37100 41076 37156 41086
rect 37100 40982 37156 41020
rect 37100 39844 37156 39854
rect 36988 39842 37156 39844
rect 36988 39790 37102 39842
rect 37154 39790 37156 39842
rect 36988 39788 37156 39790
rect 37100 39778 37156 39788
rect 36428 39554 36484 39564
rect 37100 39620 37156 39630
rect 36204 39506 36260 39518
rect 36204 39454 36206 39506
rect 36258 39454 36260 39506
rect 36204 39284 36260 39454
rect 37100 39506 37156 39564
rect 37100 39454 37102 39506
rect 37154 39454 37156 39506
rect 37100 39442 37156 39454
rect 37212 39506 37268 39518
rect 37212 39454 37214 39506
rect 37266 39454 37268 39506
rect 36316 39396 36372 39406
rect 36316 39394 36484 39396
rect 36316 39342 36318 39394
rect 36370 39342 36484 39394
rect 36316 39340 36484 39342
rect 36316 39330 36372 39340
rect 36204 39218 36260 39228
rect 34860 39006 34862 39058
rect 34914 39006 34916 39058
rect 33628 38722 33684 38734
rect 33628 38670 33630 38722
rect 33682 38670 33684 38722
rect 33628 38668 33684 38670
rect 32284 37998 32286 38050
rect 32338 37998 32340 38050
rect 32284 37986 32340 37998
rect 32956 38612 33684 38668
rect 32060 37886 32062 37938
rect 32114 37886 32116 37938
rect 32060 37874 32116 37886
rect 31948 37426 32004 37436
rect 32956 37826 33012 38612
rect 33628 38052 33684 38062
rect 33628 38050 33796 38052
rect 33628 37998 33630 38050
rect 33682 37998 33796 38050
rect 33628 37996 33796 37998
rect 33628 37986 33684 37996
rect 32956 37774 32958 37826
rect 33010 37774 33012 37826
rect 32956 37044 33012 37774
rect 32508 36988 33012 37044
rect 33740 37156 33796 37996
rect 34300 37940 34356 37950
rect 34300 37846 34356 37884
rect 30940 36372 30996 36382
rect 30940 36370 31108 36372
rect 30940 36318 30942 36370
rect 30994 36318 31108 36370
rect 30940 36316 31108 36318
rect 30940 36306 30996 36316
rect 30604 34132 30660 34142
rect 30604 34130 30772 34132
rect 30604 34078 30606 34130
rect 30658 34078 30772 34130
rect 30604 34076 30772 34078
rect 30604 34066 30660 34076
rect 30492 33292 30660 33348
rect 30268 33282 30324 33292
rect 29596 33124 29652 33134
rect 29596 32452 29652 33068
rect 30268 33122 30324 33134
rect 30268 33070 30270 33122
rect 30322 33070 30324 33122
rect 29932 32452 29988 32462
rect 29596 32450 29988 32452
rect 29596 32398 29934 32450
rect 29986 32398 29988 32450
rect 29596 32396 29988 32398
rect 29260 31892 29316 32060
rect 29932 32004 29988 32396
rect 30268 32340 30324 33070
rect 30492 33124 30548 33134
rect 30492 33030 30548 33068
rect 30380 32676 30436 32686
rect 30380 32582 30436 32620
rect 30492 32564 30548 32574
rect 30492 32470 30548 32508
rect 30380 32340 30436 32350
rect 30268 32338 30436 32340
rect 30268 32286 30382 32338
rect 30434 32286 30436 32338
rect 30268 32284 30436 32286
rect 30380 32274 30436 32284
rect 29932 31938 29988 31948
rect 29260 31890 29428 31892
rect 29260 31838 29262 31890
rect 29314 31838 29428 31890
rect 29260 31836 29428 31838
rect 29260 31826 29316 31836
rect 29372 30994 29428 31836
rect 29372 30942 29374 30994
rect 29426 30942 29428 30994
rect 29372 30930 29428 30942
rect 30156 30882 30212 30894
rect 30156 30830 30158 30882
rect 30210 30830 30212 30882
rect 30156 30548 30212 30830
rect 30156 30482 30212 30492
rect 30604 30436 30660 33292
rect 30716 33346 30772 34076
rect 30940 34018 30996 34030
rect 30940 33966 30942 34018
rect 30994 33966 30996 34018
rect 30940 33908 30996 33966
rect 30940 33842 30996 33852
rect 31052 33458 31108 36316
rect 32172 35028 32228 35038
rect 32172 34934 32228 34972
rect 31052 33406 31054 33458
rect 31106 33406 31108 33458
rect 31052 33394 31108 33406
rect 30716 33294 30718 33346
rect 30770 33294 30772 33346
rect 30716 33282 30772 33294
rect 31052 33122 31108 33134
rect 31052 33070 31054 33122
rect 31106 33070 31108 33122
rect 31052 32788 31108 33070
rect 31276 33124 31332 33134
rect 31164 32788 31220 32798
rect 31052 32786 31220 32788
rect 31052 32734 31166 32786
rect 31218 32734 31220 32786
rect 31052 32732 31220 32734
rect 31164 32722 31220 32732
rect 30940 32674 30996 32686
rect 30940 32622 30942 32674
rect 30994 32622 30996 32674
rect 30828 32564 30884 32574
rect 30828 31220 30884 32508
rect 30940 32452 30996 32622
rect 30940 32386 30996 32396
rect 31276 31892 31332 33068
rect 31500 32676 31556 32686
rect 31500 32452 31556 32620
rect 32396 32674 32452 32686
rect 32396 32622 32398 32674
rect 32450 32622 32452 32674
rect 32284 32564 32340 32574
rect 32284 32470 32340 32508
rect 31948 32452 32004 32462
rect 31500 32450 31668 32452
rect 31500 32398 31502 32450
rect 31554 32398 31668 32450
rect 31500 32396 31668 32398
rect 31500 32386 31556 32396
rect 31276 31836 31556 31892
rect 30828 31164 31332 31220
rect 30716 30548 30772 30558
rect 30772 30492 30884 30548
rect 30716 30482 30772 30492
rect 30492 30380 30660 30436
rect 30828 30434 30884 30492
rect 30828 30382 30830 30434
rect 30882 30382 30884 30434
rect 30492 30324 30548 30380
rect 30828 30370 30884 30382
rect 30380 30268 30548 30324
rect 29372 30212 29428 30222
rect 29372 30118 29428 30156
rect 29820 30212 29876 30222
rect 29708 30098 29764 30110
rect 29708 30046 29710 30098
rect 29762 30046 29764 30098
rect 29708 29540 29764 30046
rect 29820 30098 29876 30156
rect 29820 30046 29822 30098
rect 29874 30046 29876 30098
rect 29820 30034 29876 30046
rect 30044 30100 30100 30110
rect 30268 30100 30324 30110
rect 30044 30098 30324 30100
rect 30044 30046 30046 30098
rect 30098 30046 30270 30098
rect 30322 30046 30324 30098
rect 30044 30044 30324 30046
rect 30044 30034 30100 30044
rect 30268 30034 30324 30044
rect 29708 29484 30100 29540
rect 29036 28466 29092 28476
rect 29148 29426 29204 29438
rect 29148 29374 29150 29426
rect 29202 29374 29204 29426
rect 29148 29316 29204 29374
rect 29708 29316 29764 29326
rect 29148 29314 29764 29316
rect 29148 29262 29710 29314
rect 29762 29262 29764 29314
rect 29148 29260 29764 29262
rect 29148 26628 29204 29260
rect 29708 29250 29764 29260
rect 29372 28868 29428 28878
rect 30044 28868 30100 29484
rect 30380 28980 30436 30268
rect 30940 30212 30996 30222
rect 30492 30210 30996 30212
rect 30492 30158 30942 30210
rect 30994 30158 30996 30210
rect 30492 30156 30996 30158
rect 30492 30098 30548 30156
rect 30940 30146 30996 30156
rect 30492 30046 30494 30098
rect 30546 30046 30548 30098
rect 30492 30034 30548 30046
rect 31164 30100 31220 30110
rect 30716 29988 30772 29998
rect 30716 29894 30772 29932
rect 31164 29986 31220 30044
rect 31276 30100 31332 31164
rect 31276 30098 31444 30100
rect 31276 30046 31278 30098
rect 31330 30046 31444 30098
rect 31276 30044 31444 30046
rect 31276 30034 31332 30044
rect 31164 29934 31166 29986
rect 31218 29934 31220 29986
rect 30044 28812 30324 28868
rect 29372 28774 29428 28812
rect 29932 28644 29988 28654
rect 30156 28644 30212 28654
rect 29932 28642 30212 28644
rect 29932 28590 29934 28642
rect 29986 28590 30158 28642
rect 30210 28590 30212 28642
rect 29932 28588 30212 28590
rect 29932 28578 29988 28588
rect 30156 28578 30212 28588
rect 30268 28532 30324 28812
rect 30268 28466 30324 28476
rect 30380 28530 30436 28924
rect 31164 29092 31220 29934
rect 30380 28478 30382 28530
rect 30434 28478 30436 28530
rect 29484 28420 29540 28430
rect 29484 28326 29540 28364
rect 29708 28420 29764 28430
rect 30044 28420 30100 28430
rect 29708 28418 29876 28420
rect 29708 28366 29710 28418
rect 29762 28366 29876 28418
rect 29708 28364 29876 28366
rect 29708 28354 29764 28364
rect 29708 27412 29764 27422
rect 29260 27300 29316 27310
rect 29260 27298 29540 27300
rect 29260 27246 29262 27298
rect 29314 27246 29540 27298
rect 29260 27244 29540 27246
rect 29260 27234 29316 27244
rect 29372 27074 29428 27086
rect 29372 27022 29374 27074
rect 29426 27022 29428 27074
rect 29260 26964 29316 27002
rect 29260 26898 29316 26908
rect 29372 26852 29428 27022
rect 29372 26786 29428 26796
rect 29260 26628 29316 26638
rect 29148 26572 29260 26628
rect 28924 26338 28980 26348
rect 28812 26238 28814 26290
rect 28866 26238 28868 26290
rect 28812 26226 28868 26238
rect 29260 25618 29316 26572
rect 29372 26404 29428 26414
rect 29484 26404 29540 27244
rect 29708 26964 29764 27356
rect 29820 27298 29876 28364
rect 29820 27246 29822 27298
rect 29874 27246 29876 27298
rect 29820 27234 29876 27246
rect 29932 27074 29988 27086
rect 29932 27022 29934 27074
rect 29986 27022 29988 27074
rect 29820 26964 29876 26974
rect 29708 26962 29876 26964
rect 29708 26910 29822 26962
rect 29874 26910 29876 26962
rect 29708 26908 29876 26910
rect 29708 26740 29764 26908
rect 29820 26898 29876 26908
rect 29932 26852 29988 27022
rect 29932 26786 29988 26796
rect 30044 26964 30100 28364
rect 30380 28420 30436 28478
rect 30492 28642 30548 28654
rect 30492 28590 30494 28642
rect 30546 28590 30548 28642
rect 30492 28532 30548 28590
rect 30604 28532 30660 28542
rect 30492 28476 30604 28532
rect 30604 28466 30660 28476
rect 31052 28532 31108 28542
rect 30380 28354 30436 28364
rect 30940 28420 30996 28430
rect 30940 28326 30996 28364
rect 31052 28196 31108 28476
rect 30940 28140 31108 28196
rect 30604 27188 30660 27198
rect 30604 27094 30660 27132
rect 30940 27076 30996 28140
rect 31164 28084 31220 29036
rect 31388 28530 31444 30044
rect 31500 29988 31556 31836
rect 31500 29922 31556 29932
rect 31388 28478 31390 28530
rect 31442 28478 31444 28530
rect 31388 28466 31444 28478
rect 30268 26964 30324 27002
rect 30044 26908 30268 26964
rect 30716 26962 30772 26974
rect 30716 26910 30718 26962
rect 30770 26910 30772 26962
rect 30716 26908 30772 26910
rect 29708 26674 29764 26684
rect 30044 26628 30100 26908
rect 30268 26898 30324 26908
rect 30492 26850 30548 26862
rect 30492 26798 30494 26850
rect 30546 26798 30548 26850
rect 29820 26572 30100 26628
rect 30268 26740 30324 26750
rect 29820 26514 29876 26572
rect 29820 26462 29822 26514
rect 29874 26462 29876 26514
rect 29820 26450 29876 26462
rect 30268 26514 30324 26684
rect 30268 26462 30270 26514
rect 30322 26462 30324 26514
rect 29372 26402 29540 26404
rect 29372 26350 29374 26402
rect 29426 26350 29540 26402
rect 29372 26348 29540 26350
rect 29372 26338 29428 26348
rect 29596 26292 29652 26302
rect 29596 26290 29764 26292
rect 29596 26238 29598 26290
rect 29650 26238 29764 26290
rect 29596 26236 29764 26238
rect 29596 26226 29652 26236
rect 29484 26180 29540 26190
rect 29484 26086 29540 26124
rect 29708 25730 29764 26236
rect 30268 26180 30324 26462
rect 30268 26114 30324 26124
rect 30492 26068 30548 26798
rect 30604 26852 30772 26908
rect 30604 26514 30660 26852
rect 30604 26462 30606 26514
rect 30658 26462 30660 26514
rect 30604 26450 30660 26462
rect 30828 26404 30884 26414
rect 30828 26310 30884 26348
rect 30940 26402 30996 27020
rect 30940 26350 30942 26402
rect 30994 26350 30996 26402
rect 30940 26338 30996 26350
rect 31052 28028 31220 28084
rect 31052 26180 31108 28028
rect 31164 27074 31220 27086
rect 31164 27022 31166 27074
rect 31218 27022 31220 27074
rect 31164 26628 31220 27022
rect 31164 26562 31220 26572
rect 31500 26740 31556 26750
rect 31500 26404 31556 26684
rect 31500 26310 31556 26348
rect 30940 26124 31108 26180
rect 30492 26012 30884 26068
rect 29708 25678 29710 25730
rect 29762 25678 29764 25730
rect 29708 25666 29764 25678
rect 29260 25566 29262 25618
rect 29314 25566 29316 25618
rect 29260 25554 29316 25566
rect 30044 25508 30100 25518
rect 29932 25452 30044 25508
rect 29820 25396 29876 25406
rect 29820 25302 29876 25340
rect 28476 25116 28756 25172
rect 29708 25282 29764 25294
rect 29708 25230 29710 25282
rect 29762 25230 29764 25282
rect 29708 25172 29764 25230
rect 26796 24948 26852 24958
rect 26796 24612 26852 24892
rect 26796 24556 26964 24612
rect 26460 22482 26628 22484
rect 26460 22430 26462 22482
rect 26514 22430 26628 22482
rect 26460 22428 26628 22430
rect 26460 22418 26516 22428
rect 26460 22260 26516 22270
rect 26236 18398 26238 18450
rect 26290 18398 26292 18450
rect 25116 16658 25172 17164
rect 25452 17108 25508 17500
rect 25116 16606 25118 16658
rect 25170 16606 25172 16658
rect 25116 16594 25172 16606
rect 25228 17052 25508 17108
rect 25900 18340 25956 18350
rect 26236 18340 26292 18398
rect 25900 18338 26292 18340
rect 25900 18286 25902 18338
rect 25954 18286 26292 18338
rect 25900 18284 26292 18286
rect 26348 21924 26404 21934
rect 25900 17668 25956 18284
rect 26348 18228 26404 21868
rect 24108 15026 24164 15036
rect 24332 15092 24500 15148
rect 24332 13636 24388 15092
rect 25228 14420 25284 17052
rect 25340 16770 25396 16782
rect 25340 16718 25342 16770
rect 25394 16718 25396 16770
rect 25340 16658 25396 16718
rect 25340 16606 25342 16658
rect 25394 16606 25396 16658
rect 25340 15538 25396 16606
rect 25564 16772 25620 16782
rect 25564 16210 25620 16716
rect 25900 16660 25956 17612
rect 26236 18172 26404 18228
rect 25956 16604 26068 16660
rect 25900 16594 25956 16604
rect 25564 16158 25566 16210
rect 25618 16158 25620 16210
rect 25564 16146 25620 16158
rect 26012 16210 26068 16604
rect 26012 16158 26014 16210
rect 26066 16158 26068 16210
rect 26012 16146 26068 16158
rect 25340 15486 25342 15538
rect 25394 15486 25396 15538
rect 25340 15316 25396 15486
rect 25340 15250 25396 15260
rect 26236 15148 26292 18172
rect 26460 18116 26516 22204
rect 26572 22148 26628 22428
rect 26684 23714 26740 23726
rect 26684 23662 26686 23714
rect 26738 23662 26740 23714
rect 26684 23492 26740 23662
rect 26684 22484 26740 23436
rect 26908 22932 26964 24556
rect 28476 24052 28532 25116
rect 29708 25106 29764 25116
rect 29036 25060 29092 25070
rect 27916 24050 28532 24052
rect 27916 23998 28478 24050
rect 28530 23998 28532 24050
rect 27916 23996 28532 23998
rect 27916 23826 27972 23996
rect 28476 23986 28532 23996
rect 28588 24892 28980 24948
rect 27916 23774 27918 23826
rect 27970 23774 27972 23826
rect 27916 23762 27972 23774
rect 28028 23826 28084 23838
rect 28028 23774 28030 23826
rect 28082 23774 28084 23826
rect 27692 23716 27748 23726
rect 27692 23714 27860 23716
rect 27692 23662 27694 23714
rect 27746 23662 27860 23714
rect 27692 23660 27860 23662
rect 27692 23650 27748 23660
rect 27804 23156 27860 23660
rect 28028 23380 28084 23774
rect 28084 23324 28196 23380
rect 28028 23314 28084 23324
rect 27804 23100 27972 23156
rect 27244 23044 27300 23054
rect 27244 23042 27524 23044
rect 27244 22990 27246 23042
rect 27298 22990 27524 23042
rect 27244 22988 27524 22990
rect 27244 22978 27300 22988
rect 26908 22866 26964 22876
rect 27468 22596 27524 22988
rect 27468 22540 27860 22596
rect 26684 22418 26740 22428
rect 27692 22258 27748 22270
rect 27692 22206 27694 22258
rect 27746 22206 27748 22258
rect 26572 22082 26628 22092
rect 26908 22146 26964 22158
rect 26908 22094 26910 22146
rect 26962 22094 26964 22146
rect 26908 22036 26964 22094
rect 26012 15092 26292 15148
rect 26348 18060 26516 18116
rect 26684 21980 26908 22036
rect 25340 14530 25396 14542
rect 25340 14478 25342 14530
rect 25394 14478 25396 14530
rect 25340 14420 25396 14478
rect 25788 14420 25844 14430
rect 25228 14418 25844 14420
rect 25228 14366 25790 14418
rect 25842 14366 25844 14418
rect 25228 14364 25844 14366
rect 25788 14354 25844 14364
rect 24220 13634 24388 13636
rect 24220 13582 24334 13634
rect 24386 13582 24388 13634
rect 24220 13580 24388 13582
rect 24220 13076 24276 13580
rect 24332 13570 24388 13580
rect 25116 14306 25172 14318
rect 25116 14254 25118 14306
rect 25170 14254 25172 14306
rect 24780 13076 24836 13086
rect 24220 13074 24836 13076
rect 24220 13022 24782 13074
rect 24834 13022 24836 13074
rect 24220 13020 24836 13022
rect 23996 12852 24052 12862
rect 23996 12758 24052 12796
rect 24220 12850 24276 13020
rect 24780 13010 24836 13020
rect 24220 12798 24222 12850
rect 24274 12798 24276 12850
rect 24220 12786 24276 12798
rect 24332 12850 24388 12862
rect 24332 12798 24334 12850
rect 24386 12798 24388 12850
rect 24332 12628 24388 12798
rect 23884 12572 24164 12628
rect 24108 12402 24164 12572
rect 24108 12350 24110 12402
rect 24162 12350 24164 12402
rect 23884 12180 23940 12190
rect 23884 12086 23940 12124
rect 24108 11956 24164 12350
rect 24220 12572 24388 12628
rect 24220 12180 24276 12572
rect 24220 12086 24276 12124
rect 25116 12180 25172 14254
rect 25340 13636 25396 13646
rect 25228 13412 25284 13422
rect 25228 12404 25284 13356
rect 25228 12338 25284 12348
rect 25340 12740 25396 13580
rect 25676 12962 25732 12974
rect 25676 12910 25678 12962
rect 25730 12910 25732 12962
rect 25676 12740 25732 12910
rect 25340 12738 25732 12740
rect 25340 12686 25342 12738
rect 25394 12686 25732 12738
rect 25340 12684 25732 12686
rect 25116 12114 25172 12124
rect 24668 12066 24724 12078
rect 24668 12014 24670 12066
rect 24722 12014 24724 12066
rect 24668 11956 24724 12014
rect 24108 11900 24724 11956
rect 24332 11506 24388 11900
rect 24332 11454 24334 11506
rect 24386 11454 24388 11506
rect 24332 11442 24388 11454
rect 23100 9774 23102 9826
rect 23154 9774 23156 9826
rect 23100 9762 23156 9774
rect 24780 11172 24836 11182
rect 21420 9604 21476 9614
rect 20972 8418 21028 8428
rect 21308 9602 21476 9604
rect 21308 9550 21422 9602
rect 21474 9550 21476 9602
rect 21308 9548 21476 9550
rect 20524 8260 20580 8270
rect 20524 8166 20580 8204
rect 20748 8258 20804 8270
rect 20748 8206 20750 8258
rect 20802 8206 20804 8258
rect 20412 8148 20468 8158
rect 20412 8054 20468 8092
rect 19628 7494 19684 7532
rect 19740 7698 20244 7700
rect 19740 7646 20078 7698
rect 20130 7646 20244 7698
rect 19740 7644 20244 7646
rect 20300 8034 20356 8046
rect 20300 7982 20302 8034
rect 20354 7982 20356 8034
rect 20300 7924 20356 7982
rect 20748 8036 20804 8206
rect 20748 7970 20804 7980
rect 18284 6750 18286 6802
rect 18338 6750 18340 6802
rect 18284 6738 18340 6750
rect 19516 7476 19572 7486
rect 16156 6638 16158 6690
rect 16210 6638 16212 6690
rect 16156 6626 16212 6638
rect 14700 6078 14702 6130
rect 14754 6078 14756 6130
rect 14588 5124 14644 5134
rect 14700 5124 14756 6078
rect 19516 6132 19572 7420
rect 19740 7364 19796 7644
rect 20076 7634 20132 7644
rect 19852 7476 19908 7486
rect 19852 7382 19908 7420
rect 20188 7474 20244 7486
rect 20188 7422 20190 7474
rect 20242 7422 20244 7474
rect 19516 6066 19572 6076
rect 19628 7308 19796 7364
rect 19964 7364 20020 7374
rect 18956 6018 19012 6030
rect 18956 5966 18958 6018
rect 19010 5966 19012 6018
rect 17388 5908 17444 5918
rect 15260 5684 15316 5694
rect 15260 5234 15316 5628
rect 15260 5182 15262 5234
rect 15314 5182 15316 5234
rect 15260 5170 15316 5182
rect 17388 5234 17444 5852
rect 18844 5684 18900 5694
rect 18844 5590 18900 5628
rect 18844 5236 18900 5246
rect 17388 5182 17390 5234
rect 17442 5182 17444 5234
rect 17388 5170 17444 5182
rect 18172 5234 18900 5236
rect 18172 5182 18846 5234
rect 18898 5182 18900 5234
rect 18172 5180 18900 5182
rect 14588 5122 14700 5124
rect 14588 5070 14590 5122
rect 14642 5070 14700 5122
rect 14588 5068 14700 5070
rect 14588 5058 14644 5068
rect 14700 5030 14756 5068
rect 16828 5124 16884 5134
rect 16828 4564 16884 5068
rect 17836 5124 17892 5134
rect 17836 5030 17892 5068
rect 16828 4562 17444 4564
rect 16828 4510 16830 4562
rect 16882 4510 17444 4562
rect 16828 4508 17444 4510
rect 16828 4498 16884 4508
rect 14364 4452 14420 4462
rect 14364 4338 14420 4396
rect 14924 4452 14980 4462
rect 14924 4358 14980 4396
rect 14364 4286 14366 4338
rect 14418 4286 14420 4338
rect 14364 4274 14420 4286
rect 17388 4338 17444 4508
rect 18172 4450 18228 5180
rect 18844 5170 18900 5180
rect 18956 5124 19012 5966
rect 19628 5908 19684 7308
rect 19964 7270 20020 7308
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19740 6132 19796 6142
rect 19740 6038 19796 6076
rect 20188 6132 20244 7422
rect 20300 7476 20356 7868
rect 20860 7700 20916 7710
rect 20860 7606 20916 7644
rect 20300 7410 20356 7420
rect 20636 7364 20692 7374
rect 20636 7270 20692 7308
rect 20748 7362 20804 7374
rect 20748 7310 20750 7362
rect 20802 7310 20804 7362
rect 20748 6804 20804 7310
rect 20748 6738 20804 6748
rect 19964 6020 20020 6030
rect 19964 5926 20020 5964
rect 19628 5814 19684 5852
rect 20188 5906 20244 6076
rect 20188 5854 20190 5906
rect 20242 5854 20244 5906
rect 20188 5842 20244 5854
rect 20300 6020 20356 6030
rect 19852 5794 19908 5806
rect 19852 5742 19854 5794
rect 19906 5742 19908 5794
rect 19180 5684 19236 5694
rect 19852 5684 19908 5742
rect 19180 5682 19908 5684
rect 19180 5630 19182 5682
rect 19234 5630 19908 5682
rect 19180 5628 19908 5630
rect 19180 5618 19236 5628
rect 19180 5348 19236 5358
rect 19180 5254 19236 5292
rect 18956 5010 19012 5068
rect 18956 4958 18958 5010
rect 19010 4958 19012 5010
rect 18956 4946 19012 4958
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 18172 4398 18174 4450
rect 18226 4398 18228 4450
rect 18172 4386 18228 4398
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 17388 4274 17444 4286
rect 20300 4226 20356 5964
rect 21308 6020 21364 9548
rect 21420 9538 21476 9548
rect 21980 9602 22036 9614
rect 22876 9604 22932 9614
rect 21980 9550 21982 9602
rect 22034 9550 22036 9602
rect 21980 8260 22036 9550
rect 21980 8194 22036 8204
rect 22204 9602 22932 9604
rect 22204 9550 22878 9602
rect 22930 9550 22932 9602
rect 22204 9548 22932 9550
rect 22204 8932 22260 9548
rect 22876 9538 22932 9548
rect 22204 8258 22260 8876
rect 22204 8206 22206 8258
rect 22258 8206 22260 8258
rect 22204 8194 22260 8206
rect 22652 8260 22708 8270
rect 22652 8166 22708 8204
rect 23100 8258 23156 8270
rect 23100 8206 23102 8258
rect 23154 8206 23156 8258
rect 22092 8036 22148 8046
rect 21980 7586 22036 7598
rect 21980 7534 21982 7586
rect 22034 7534 22036 7586
rect 21644 6468 21700 6478
rect 21644 6130 21700 6412
rect 21644 6078 21646 6130
rect 21698 6078 21700 6130
rect 21644 6066 21700 6078
rect 21756 6132 21812 6142
rect 21980 6132 22036 7534
rect 22092 7476 22148 7980
rect 22316 8034 22372 8046
rect 22316 7982 22318 8034
rect 22370 7982 22372 8034
rect 22316 7700 22372 7982
rect 22428 8034 22484 8046
rect 22428 7982 22430 8034
rect 22482 7982 22484 8034
rect 22428 7924 22484 7982
rect 23100 8036 23156 8206
rect 23772 8148 23828 8158
rect 23100 7970 23156 7980
rect 23660 8146 23828 8148
rect 23660 8094 23774 8146
rect 23826 8094 23828 8146
rect 23660 8092 23828 8094
rect 22428 7858 22484 7868
rect 23548 7700 23604 7710
rect 22316 7644 23380 7700
rect 23324 7586 23380 7644
rect 23324 7534 23326 7586
rect 23378 7534 23380 7586
rect 23324 7522 23380 7534
rect 22316 7476 22372 7486
rect 22092 7420 22316 7476
rect 22316 7382 22372 7420
rect 23548 7140 23604 7644
rect 23660 7362 23716 8092
rect 23772 8082 23828 8092
rect 24780 8036 24836 11116
rect 25340 11172 25396 12684
rect 25564 12404 25620 12414
rect 25564 11788 25620 12348
rect 25340 11106 25396 11116
rect 25452 11732 25620 11788
rect 25228 10722 25284 10734
rect 25228 10670 25230 10722
rect 25282 10670 25284 10722
rect 25228 10276 25284 10670
rect 25116 10220 25284 10276
rect 25116 9940 25172 10220
rect 25116 9874 25172 9884
rect 25340 9268 25396 9278
rect 25452 9268 25508 11732
rect 26012 11396 26068 15092
rect 26124 14308 26180 14318
rect 26124 14214 26180 14252
rect 26348 13412 26404 18060
rect 26460 15202 26516 15214
rect 26460 15150 26462 15202
rect 26514 15150 26516 15202
rect 26460 13636 26516 15150
rect 26572 14308 26628 14318
rect 26572 14214 26628 14252
rect 26460 13570 26516 13580
rect 26348 13346 26404 13356
rect 26684 13076 26740 21980
rect 26908 21970 26964 21980
rect 27020 21700 27076 21710
rect 27020 20804 27076 21644
rect 27692 21700 27748 22206
rect 27804 22148 27860 22540
rect 27916 22370 27972 23100
rect 27916 22318 27918 22370
rect 27970 22318 27972 22370
rect 27916 22306 27972 22318
rect 28028 22148 28084 22158
rect 27804 22146 28084 22148
rect 27804 22094 28030 22146
rect 28082 22094 28084 22146
rect 27804 22092 28084 22094
rect 28028 22082 28084 22092
rect 28140 21924 28196 23324
rect 28252 22372 28308 22382
rect 28252 22278 28308 22316
rect 27692 21634 27748 21644
rect 28028 21868 28196 21924
rect 27020 20710 27076 20748
rect 27692 20802 27748 20814
rect 27692 20750 27694 20802
rect 27746 20750 27748 20802
rect 27244 20690 27300 20702
rect 27244 20638 27246 20690
rect 27298 20638 27300 20690
rect 27244 20132 27300 20638
rect 27692 20692 27748 20750
rect 27916 20804 27972 20814
rect 27916 20710 27972 20748
rect 27692 20626 27748 20636
rect 27244 20066 27300 20076
rect 27356 20578 27412 20590
rect 27356 20526 27358 20578
rect 27410 20526 27412 20578
rect 27356 19236 27412 20526
rect 27916 20468 27972 20478
rect 27916 20188 27972 20412
rect 27020 19180 27412 19236
rect 27580 20132 27972 20188
rect 27020 18450 27076 19180
rect 27020 18398 27022 18450
rect 27074 18398 27076 18450
rect 27020 18386 27076 18398
rect 27580 15426 27636 20132
rect 28028 20020 28084 21868
rect 28252 20802 28308 20814
rect 28252 20750 28254 20802
rect 28306 20750 28308 20802
rect 28252 20244 28308 20750
rect 28476 20804 28532 20814
rect 28476 20710 28532 20748
rect 28364 20578 28420 20590
rect 28364 20526 28366 20578
rect 28418 20526 28420 20578
rect 28364 20468 28420 20526
rect 28364 20402 28420 20412
rect 28364 20244 28420 20254
rect 28252 20242 28420 20244
rect 28252 20190 28366 20242
rect 28418 20190 28420 20242
rect 28252 20188 28420 20190
rect 28364 20178 28420 20188
rect 28476 20242 28532 20254
rect 28476 20190 28478 20242
rect 28530 20190 28532 20242
rect 28028 19926 28084 19964
rect 28140 20130 28196 20142
rect 28140 20078 28142 20130
rect 28194 20078 28196 20130
rect 27580 15374 27582 15426
rect 27634 15374 27636 15426
rect 27580 15362 27636 15374
rect 27692 19906 27748 19918
rect 27692 19854 27694 19906
rect 27746 19854 27748 19906
rect 27692 19796 27748 19854
rect 28140 19908 28196 20078
rect 28476 20132 28532 20190
rect 28476 20066 28532 20076
rect 28140 19796 28196 19852
rect 27692 19740 28196 19796
rect 26796 15314 26852 15326
rect 26796 15262 26798 15314
rect 26850 15262 26852 15314
rect 26796 13636 26852 15262
rect 27132 13746 27188 13758
rect 27132 13694 27134 13746
rect 27186 13694 27188 13746
rect 27132 13636 27188 13694
rect 27692 13748 27748 19740
rect 27916 14308 27972 14318
rect 27916 13858 27972 14252
rect 27916 13806 27918 13858
rect 27970 13806 27972 13858
rect 27916 13794 27972 13806
rect 27692 13682 27748 13692
rect 26852 13580 27188 13636
rect 26796 13542 26852 13580
rect 26684 13010 26740 13020
rect 26460 12852 26516 12862
rect 26460 12850 27076 12852
rect 26460 12798 26462 12850
rect 26514 12798 27076 12850
rect 26460 12796 27076 12798
rect 26460 12786 26516 12796
rect 27020 12402 27076 12796
rect 27020 12350 27022 12402
rect 27074 12350 27076 12402
rect 27020 12338 27076 12350
rect 27132 12404 27188 13580
rect 27692 13076 27748 13086
rect 27132 12338 27188 12348
rect 27244 12348 27636 12404
rect 26684 12178 26740 12190
rect 26908 12180 26964 12190
rect 26684 12126 26686 12178
rect 26738 12126 26740 12178
rect 26012 11394 26180 11396
rect 26012 11342 26014 11394
rect 26066 11342 26180 11394
rect 26012 11340 26180 11342
rect 26012 11330 26068 11340
rect 25564 10610 25620 10622
rect 25564 10558 25566 10610
rect 25618 10558 25620 10610
rect 25564 9940 25620 10558
rect 26012 10498 26068 10510
rect 26012 10446 26014 10498
rect 26066 10446 26068 10498
rect 25788 9940 25844 9950
rect 26012 9940 26068 10446
rect 25564 9884 25788 9940
rect 25844 9884 26068 9940
rect 25788 9826 25844 9884
rect 25788 9774 25790 9826
rect 25842 9774 25844 9826
rect 25788 9762 25844 9774
rect 25340 9266 25508 9268
rect 25340 9214 25342 9266
rect 25394 9214 25508 9266
rect 25340 9212 25508 9214
rect 26012 9602 26068 9614
rect 26012 9550 26014 9602
rect 26066 9550 26068 9602
rect 25340 9202 25396 9212
rect 25564 9154 25620 9166
rect 25564 9102 25566 9154
rect 25618 9102 25620 9154
rect 25564 8260 25620 9102
rect 25564 8194 25620 8204
rect 25676 9044 25732 9054
rect 26012 9044 26068 9550
rect 25676 9042 26068 9044
rect 25676 8990 25678 9042
rect 25730 8990 26068 9042
rect 25676 8988 26068 8990
rect 24780 7970 24836 7980
rect 25676 7588 25732 8988
rect 25900 8370 25956 8382
rect 25900 8318 25902 8370
rect 25954 8318 25956 8370
rect 25900 8260 25956 8318
rect 25900 8194 25956 8204
rect 25676 7522 25732 7532
rect 26124 7364 26180 11340
rect 26236 11284 26292 11294
rect 26236 11190 26292 11228
rect 26684 11284 26740 12126
rect 26684 11218 26740 11228
rect 26796 12178 26964 12180
rect 26796 12126 26910 12178
rect 26962 12126 26964 12178
rect 26796 12124 26964 12126
rect 26460 9940 26516 9950
rect 26460 9846 26516 9884
rect 26572 8930 26628 8942
rect 26572 8878 26574 8930
rect 26626 8878 26628 8930
rect 26572 8484 26628 8878
rect 26572 8418 26628 8428
rect 23660 7310 23662 7362
rect 23714 7310 23716 7362
rect 23660 7298 23716 7310
rect 25564 7308 26180 7364
rect 26348 8036 26404 8046
rect 23548 7074 23604 7084
rect 25564 6690 25620 7308
rect 25564 6638 25566 6690
rect 25618 6638 25620 6690
rect 22876 6468 22932 6478
rect 22428 6244 22484 6254
rect 21812 6076 22260 6132
rect 21756 6038 21812 6076
rect 21308 5906 21364 5964
rect 21308 5854 21310 5906
rect 21362 5854 21364 5906
rect 21308 5842 21364 5854
rect 21420 5908 21476 5918
rect 21420 5814 21476 5852
rect 22204 5906 22260 6076
rect 22428 6130 22484 6188
rect 22428 6078 22430 6130
rect 22482 6078 22484 6130
rect 22428 6066 22484 6078
rect 22876 6018 22932 6412
rect 22876 5966 22878 6018
rect 22930 5966 22932 6018
rect 22876 5954 22932 5966
rect 24444 6468 24500 6478
rect 22204 5854 22206 5906
rect 22258 5854 22260 5906
rect 22204 5842 22260 5854
rect 22652 5908 22708 5918
rect 22652 5814 22708 5852
rect 21532 5794 21588 5806
rect 21532 5742 21534 5794
rect 21586 5742 21588 5794
rect 21532 5348 21588 5742
rect 22540 5794 22596 5806
rect 22540 5742 22542 5794
rect 22594 5742 22596 5794
rect 22540 5348 22596 5742
rect 22764 5348 22820 5358
rect 22540 5346 22820 5348
rect 22540 5294 22766 5346
rect 22818 5294 22820 5346
rect 22540 5292 22820 5294
rect 21532 5282 21588 5292
rect 22764 5282 22820 5292
rect 22428 5234 22484 5246
rect 22428 5182 22430 5234
rect 22482 5182 22484 5234
rect 22316 4452 22372 4462
rect 22428 4452 22484 5182
rect 22540 5124 22596 5134
rect 22540 5010 22596 5068
rect 22540 4958 22542 5010
rect 22594 4958 22596 5010
rect 22540 4946 22596 4958
rect 22316 4450 22484 4452
rect 22316 4398 22318 4450
rect 22370 4398 22484 4450
rect 22316 4396 22484 4398
rect 22316 4386 22372 4396
rect 21644 4340 21700 4350
rect 21644 4246 21700 4284
rect 20300 4174 20302 4226
rect 20354 4174 20356 4226
rect 20300 4162 20356 4174
rect 24444 4226 24500 6412
rect 25564 6130 25620 6638
rect 25788 7140 25844 7150
rect 25788 6578 25844 7084
rect 25788 6526 25790 6578
rect 25842 6526 25844 6578
rect 25788 6514 25844 6526
rect 25564 6078 25566 6130
rect 25618 6078 25620 6130
rect 25564 6066 25620 6078
rect 25228 6018 25284 6030
rect 25228 5966 25230 6018
rect 25282 5966 25284 6018
rect 25228 5124 25284 5966
rect 25228 5058 25284 5068
rect 25788 5124 25844 5134
rect 25788 5030 25844 5068
rect 26124 5124 26180 5134
rect 26124 5030 26180 5068
rect 24668 4898 24724 4910
rect 24668 4846 24670 4898
rect 24722 4846 24724 4898
rect 24668 4340 24724 4846
rect 26012 4898 26068 4910
rect 26012 4846 26014 4898
rect 26066 4846 26068 4898
rect 26012 4450 26068 4846
rect 26012 4398 26014 4450
rect 26066 4398 26068 4450
rect 26012 4386 26068 4398
rect 25228 4340 25284 4350
rect 24668 4274 24724 4284
rect 25004 4284 25228 4340
rect 24444 4174 24446 4226
rect 24498 4174 24500 4226
rect 24444 4162 24500 4174
rect 12124 4116 12180 4126
rect 10780 3490 10836 3500
rect 11676 4114 12180 4116
rect 11676 4062 12126 4114
rect 12178 4062 12180 4114
rect 11676 4060 12180 4062
rect 3276 3390 3278 3442
rect 3330 3390 3332 3442
rect 3276 3378 3332 3390
rect 7196 3444 7252 3454
rect 7196 800 7252 3388
rect 10108 3444 10164 3454
rect 10108 3350 10164 3388
rect 11676 800 11732 4060
rect 12124 4050 12180 4060
rect 11900 3668 11956 3678
rect 11900 3554 11956 3612
rect 12460 3668 12516 3678
rect 12460 3574 12516 3612
rect 25004 3666 25060 4284
rect 25228 4246 25284 4284
rect 26348 4340 26404 7980
rect 26796 6914 26852 12124
rect 26908 12114 26964 12124
rect 27244 12180 27300 12348
rect 27580 12290 27636 12348
rect 27692 12402 27748 13020
rect 28588 13076 28644 24892
rect 28924 24834 28980 24892
rect 28924 24782 28926 24834
rect 28978 24782 28980 24834
rect 28924 24770 28980 24782
rect 28812 24724 28868 24734
rect 28812 24612 28868 24668
rect 29036 24612 29092 25004
rect 29148 24948 29204 24958
rect 29148 24854 29204 24892
rect 28812 24556 29092 24612
rect 29372 23044 29428 23054
rect 29148 22372 29204 22382
rect 29148 22278 29204 22316
rect 29372 22258 29428 22988
rect 29372 22206 29374 22258
rect 29426 22206 29428 22258
rect 29372 22194 29428 22206
rect 29484 22260 29540 22270
rect 29372 20804 29428 20814
rect 29484 20804 29540 22204
rect 29372 20802 29540 20804
rect 29372 20750 29374 20802
rect 29426 20750 29540 20802
rect 29372 20748 29540 20750
rect 29820 20916 29876 20926
rect 29932 20916 29988 25452
rect 30044 25442 30100 25452
rect 30828 25506 30884 26012
rect 30828 25454 30830 25506
rect 30882 25454 30884 25506
rect 30828 25442 30884 25454
rect 30380 25284 30436 25294
rect 30940 25284 30996 26124
rect 31388 25732 31444 25742
rect 30380 25190 30436 25228
rect 30716 25228 30996 25284
rect 31052 25730 31444 25732
rect 31052 25678 31390 25730
rect 31442 25678 31444 25730
rect 31052 25676 31444 25678
rect 31052 25282 31108 25676
rect 31388 25666 31444 25676
rect 31164 25396 31220 25406
rect 31164 25302 31220 25340
rect 31052 25230 31054 25282
rect 31106 25230 31108 25282
rect 29820 20914 29988 20916
rect 29820 20862 29822 20914
rect 29874 20862 29988 20914
rect 29820 20860 29988 20862
rect 30380 23044 30436 23054
rect 29372 20738 29428 20748
rect 29036 20692 29092 20702
rect 29036 20598 29092 20636
rect 29260 20580 29316 20590
rect 29820 20580 29876 20860
rect 30268 20804 30324 20814
rect 30268 20710 30324 20748
rect 29260 20578 29876 20580
rect 29260 20526 29262 20578
rect 29314 20526 29876 20578
rect 29260 20524 29876 20526
rect 29260 20514 29316 20524
rect 28700 20130 28756 20142
rect 28700 20078 28702 20130
rect 28754 20078 28756 20130
rect 28700 19684 28756 20078
rect 28812 20020 28868 20030
rect 28812 19926 28868 19964
rect 28700 19618 28756 19628
rect 29260 19906 29316 19918
rect 29260 19854 29262 19906
rect 29314 19854 29316 19906
rect 29260 19684 29316 19854
rect 29260 19618 29316 19628
rect 29260 18676 29316 18686
rect 29372 18676 29428 20524
rect 30044 20244 30100 20282
rect 29260 18674 29428 18676
rect 29260 18622 29262 18674
rect 29314 18622 29428 18674
rect 29260 18620 29428 18622
rect 29820 20132 30100 20188
rect 29260 15204 29316 18620
rect 29596 17668 29652 17678
rect 29596 17574 29652 17612
rect 29820 16212 29876 20132
rect 30380 19236 30436 22988
rect 30604 21700 30660 21710
rect 30604 20802 30660 21644
rect 30716 21588 30772 25228
rect 30940 23716 30996 23726
rect 30828 23266 30884 23278
rect 30828 23214 30830 23266
rect 30882 23214 30884 23266
rect 30828 22260 30884 23214
rect 30828 21924 30884 22204
rect 30828 21858 30884 21868
rect 30940 21700 30996 23660
rect 30940 21634 30996 21644
rect 30828 21588 30884 21598
rect 30716 21532 30828 21588
rect 30828 21522 30884 21532
rect 30604 20750 30606 20802
rect 30658 20750 30660 20802
rect 30604 20738 30660 20750
rect 30940 20802 30996 20814
rect 30940 20750 30942 20802
rect 30994 20750 30996 20802
rect 30492 20578 30548 20590
rect 30492 20526 30494 20578
rect 30546 20526 30548 20578
rect 30492 20244 30548 20526
rect 30940 20188 30996 20750
rect 30492 20178 30548 20188
rect 30604 20132 30996 20188
rect 30604 20130 30660 20132
rect 30604 20078 30606 20130
rect 30658 20078 30660 20130
rect 30492 19236 30548 19246
rect 30380 19234 30548 19236
rect 30380 19182 30494 19234
rect 30546 19182 30548 19234
rect 30380 19180 30548 19182
rect 30492 19170 30548 19180
rect 30044 17668 30100 17678
rect 30604 17668 30660 20078
rect 31052 19684 31108 25230
rect 31388 24836 31444 24846
rect 31164 24724 31220 24734
rect 31164 24630 31220 24668
rect 31388 24722 31444 24780
rect 31388 24670 31390 24722
rect 31442 24670 31444 24722
rect 31388 24658 31444 24670
rect 31276 24500 31332 24510
rect 31276 23940 31332 24444
rect 31164 23938 31332 23940
rect 31164 23886 31278 23938
rect 31330 23886 31332 23938
rect 31164 23884 31332 23886
rect 31164 23378 31220 23884
rect 31276 23874 31332 23884
rect 31612 23716 31668 32396
rect 32004 32396 32116 32452
rect 31948 32358 32004 32396
rect 31948 31556 32004 31566
rect 31948 31462 32004 31500
rect 31836 30100 31892 30110
rect 31836 30006 31892 30044
rect 31724 28418 31780 28430
rect 31724 28366 31726 28418
rect 31778 28366 31780 28418
rect 31724 26852 31780 28366
rect 31836 27972 31892 27982
rect 31836 27878 31892 27916
rect 31836 27188 31892 27198
rect 31836 27094 31892 27132
rect 31780 26796 31892 26852
rect 31724 26786 31780 26796
rect 31724 25730 31780 25742
rect 31724 25678 31726 25730
rect 31778 25678 31780 25730
rect 31724 25618 31780 25678
rect 31724 25566 31726 25618
rect 31778 25566 31780 25618
rect 31724 25554 31780 25566
rect 31836 25396 31892 26796
rect 31836 25330 31892 25340
rect 31724 24498 31780 24510
rect 31724 24446 31726 24498
rect 31778 24446 31780 24498
rect 31724 23940 31780 24446
rect 31836 23940 31892 23950
rect 31724 23938 31892 23940
rect 31724 23886 31838 23938
rect 31890 23886 31892 23938
rect 31724 23884 31892 23886
rect 31164 23326 31166 23378
rect 31218 23326 31220 23378
rect 31164 23314 31220 23326
rect 31276 23660 31668 23716
rect 30828 19346 30884 19358
rect 30828 19294 30830 19346
rect 30882 19294 30884 19346
rect 30716 19012 30772 19022
rect 30716 17778 30772 18956
rect 30716 17726 30718 17778
rect 30770 17726 30772 17778
rect 30716 17714 30772 17726
rect 30100 17612 30660 17668
rect 30044 17574 30100 17612
rect 29820 15538 29876 16156
rect 29820 15486 29822 15538
rect 29874 15486 29876 15538
rect 29820 15474 29876 15486
rect 30716 15316 30772 15326
rect 30828 15316 30884 19294
rect 30940 18900 30996 18910
rect 30940 18004 30996 18844
rect 31052 18228 31108 19628
rect 31164 19460 31220 19470
rect 31164 19346 31220 19404
rect 31164 19294 31166 19346
rect 31218 19294 31220 19346
rect 31164 19282 31220 19294
rect 31052 18162 31108 18172
rect 31164 19124 31220 19134
rect 30940 17948 31108 18004
rect 29260 15138 29316 15148
rect 30044 15314 30884 15316
rect 30044 15262 30718 15314
rect 30770 15262 30884 15314
rect 30044 15260 30884 15262
rect 30940 15426 30996 15438
rect 30940 15374 30942 15426
rect 30994 15374 30996 15426
rect 30044 13634 30100 15260
rect 30716 15250 30772 15260
rect 30940 15092 30996 15374
rect 30940 15026 30996 15036
rect 30044 13582 30046 13634
rect 30098 13582 30100 13634
rect 30044 13570 30100 13582
rect 31052 13300 31108 17948
rect 31164 13860 31220 19068
rect 31276 18900 31332 23660
rect 31500 23380 31556 23390
rect 31500 19234 31556 23324
rect 31836 23378 31892 23884
rect 31836 23326 31838 23378
rect 31890 23326 31892 23378
rect 31836 23314 31892 23326
rect 31612 21588 31668 21598
rect 31612 19908 31668 21532
rect 31724 21476 31780 21486
rect 31724 20914 31780 21420
rect 31724 20862 31726 20914
rect 31778 20862 31780 20914
rect 31724 20850 31780 20862
rect 31612 19842 31668 19852
rect 32060 20804 32116 32396
rect 32396 31556 32452 32622
rect 32508 31780 32564 36988
rect 33180 36258 33236 36270
rect 33180 36206 33182 36258
rect 33234 36206 33236 36258
rect 33068 35698 33124 35710
rect 33068 35646 33070 35698
rect 33122 35646 33124 35698
rect 32732 35364 32788 35374
rect 32732 35026 32788 35308
rect 33068 35364 33124 35646
rect 33068 35298 33124 35308
rect 32732 34974 32734 35026
rect 32786 34974 32788 35026
rect 32732 34962 32788 34974
rect 33180 34580 33236 36206
rect 33740 36258 33796 37100
rect 33740 36206 33742 36258
rect 33794 36206 33796 36258
rect 33068 34524 33236 34580
rect 33516 35364 33572 35374
rect 33740 35364 33796 36206
rect 33572 35308 33796 35364
rect 33852 35586 33908 35598
rect 33852 35534 33854 35586
rect 33906 35534 33908 35586
rect 33068 33908 33124 34524
rect 33068 33842 33124 33852
rect 33180 34356 33236 34366
rect 33180 33570 33236 34300
rect 33180 33518 33182 33570
rect 33234 33518 33236 33570
rect 33180 33506 33236 33518
rect 33516 33460 33572 35308
rect 33852 34356 33908 35534
rect 33852 34290 33908 34300
rect 33516 33404 33684 33460
rect 33180 33348 33236 33358
rect 32844 33124 32900 33134
rect 33068 33124 33124 33134
rect 32844 33030 32900 33068
rect 32956 33122 33124 33124
rect 32956 33070 33070 33122
rect 33122 33070 33124 33122
rect 32956 33068 33124 33070
rect 32620 32676 32676 32686
rect 32956 32676 33012 33068
rect 33068 33058 33124 33068
rect 33180 32788 33236 33292
rect 33292 33236 33348 33246
rect 33516 33236 33572 33246
rect 33292 33234 33572 33236
rect 33292 33182 33294 33234
rect 33346 33182 33518 33234
rect 33570 33182 33572 33234
rect 33292 33180 33572 33182
rect 33292 33170 33348 33180
rect 33516 33170 33572 33180
rect 33404 32788 33460 32798
rect 33180 32786 33460 32788
rect 33180 32734 33406 32786
rect 33458 32734 33460 32786
rect 33180 32732 33460 32734
rect 33404 32722 33460 32732
rect 32620 32674 33012 32676
rect 32620 32622 32622 32674
rect 32674 32622 33012 32674
rect 32620 32620 33012 32622
rect 32620 32610 32676 32620
rect 32508 31714 32564 31724
rect 33180 32564 33236 32574
rect 32396 31490 32452 31500
rect 33180 31218 33236 32508
rect 33516 32564 33572 32574
rect 33628 32564 33684 33404
rect 33852 33348 33908 33358
rect 33908 33292 34132 33348
rect 33852 33254 33908 33292
rect 33740 33236 33796 33246
rect 33740 33142 33796 33180
rect 34076 32786 34132 33292
rect 34300 33236 34356 33246
rect 34300 33142 34356 33180
rect 34076 32734 34078 32786
rect 34130 32734 34132 32786
rect 34076 32722 34132 32734
rect 34300 32674 34356 32686
rect 34300 32622 34302 32674
rect 34354 32622 34356 32674
rect 33572 32508 33684 32564
rect 33740 32564 33796 32574
rect 33740 32562 33908 32564
rect 33740 32510 33742 32562
rect 33794 32510 33908 32562
rect 33740 32508 33908 32510
rect 33516 32498 33572 32508
rect 33740 32498 33796 32508
rect 33740 32116 33796 32126
rect 33516 31892 33572 31902
rect 33180 31166 33182 31218
rect 33234 31166 33236 31218
rect 33180 31154 33236 31166
rect 33292 31556 33348 31566
rect 32396 30882 32452 30894
rect 32396 30830 32398 30882
rect 32450 30830 32452 30882
rect 32396 30212 32452 30830
rect 32396 29428 32452 30156
rect 32396 29362 32452 29372
rect 33292 30324 33348 31500
rect 33516 31556 33572 31836
rect 33516 31490 33572 31500
rect 33740 31554 33796 32060
rect 33740 31502 33742 31554
rect 33794 31502 33796 31554
rect 32172 28868 32228 28878
rect 32172 24946 32228 28812
rect 32172 24894 32174 24946
rect 32226 24894 32228 24946
rect 32172 24724 32228 24894
rect 32284 25172 32340 25182
rect 32284 24836 32340 25116
rect 33292 24948 33348 30268
rect 33740 30884 33796 31502
rect 33852 31332 33908 32508
rect 34300 32116 34356 32622
rect 34524 32564 34580 32574
rect 34524 32562 34692 32564
rect 34524 32510 34526 32562
rect 34578 32510 34692 32562
rect 34524 32508 34692 32510
rect 34524 32498 34580 32508
rect 34412 32452 34468 32462
rect 34412 32358 34468 32396
rect 34300 32050 34356 32060
rect 34636 32002 34692 32508
rect 34636 31950 34638 32002
rect 34690 31950 34692 32002
rect 34636 31938 34692 31950
rect 34748 32562 34804 32574
rect 34748 32510 34750 32562
rect 34802 32510 34804 32562
rect 34748 31892 34804 32510
rect 34748 31826 34804 31836
rect 34636 31610 34692 31622
rect 34636 31558 34638 31610
rect 34690 31558 34692 31610
rect 34636 31556 34692 31558
rect 34636 31490 34692 31500
rect 34748 31610 34804 31622
rect 34748 31558 34750 31610
rect 34802 31558 34804 31610
rect 34748 31332 34804 31558
rect 33852 31266 33908 31276
rect 34636 31276 34748 31332
rect 33628 29988 33684 29998
rect 33628 29894 33684 29932
rect 33740 29652 33796 30828
rect 34636 30212 34692 31276
rect 34748 31266 34804 31276
rect 34636 30118 34692 30156
rect 33964 29988 34020 29998
rect 34300 29988 34356 29998
rect 33964 29894 34020 29932
rect 34188 29986 34356 29988
rect 34188 29934 34302 29986
rect 34354 29934 34356 29986
rect 34188 29932 34356 29934
rect 33740 29586 33796 29596
rect 33964 29538 34020 29550
rect 33964 29486 33966 29538
rect 34018 29486 34020 29538
rect 33964 27524 34020 29486
rect 34188 28532 34244 29932
rect 34300 29922 34356 29932
rect 34412 29988 34468 29998
rect 34300 29652 34356 29662
rect 34412 29652 34468 29932
rect 34300 29650 34468 29652
rect 34300 29598 34302 29650
rect 34354 29598 34468 29650
rect 34300 29596 34468 29598
rect 34300 29586 34356 29596
rect 34188 28466 34244 28476
rect 34076 28420 34132 28430
rect 34076 28082 34132 28364
rect 34076 28030 34078 28082
rect 34130 28030 34132 28082
rect 34076 27972 34132 28030
rect 34748 28420 34804 28430
rect 34748 28082 34804 28364
rect 34748 28030 34750 28082
rect 34802 28030 34804 28082
rect 34748 28018 34804 28030
rect 34300 27972 34356 27982
rect 34076 27970 34356 27972
rect 34076 27918 34302 27970
rect 34354 27918 34356 27970
rect 34076 27916 34356 27918
rect 34300 27906 34356 27916
rect 34860 27972 34916 39006
rect 36316 38722 36372 38734
rect 36316 38670 36318 38722
rect 36370 38670 36372 38722
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 36316 37156 36372 38670
rect 36428 38164 36484 39340
rect 36540 39394 36596 39406
rect 36540 39342 36542 39394
rect 36594 39342 36596 39394
rect 36540 38668 36596 39342
rect 37212 39284 37268 39454
rect 37212 39218 37268 39228
rect 36540 38612 37044 38668
rect 36428 38162 36708 38164
rect 36428 38110 36430 38162
rect 36482 38110 36708 38162
rect 36428 38108 36708 38110
rect 36428 38098 36484 38108
rect 36428 37156 36484 37166
rect 36316 37100 36428 37156
rect 36428 37062 36484 37100
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 36204 36372 36260 36382
rect 36204 36278 36260 36316
rect 35756 36258 35812 36270
rect 35756 36206 35758 36258
rect 35810 36206 35812 36258
rect 35756 35924 35812 36206
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35756 35028 35812 35868
rect 36540 35810 36596 35822
rect 36540 35758 36542 35810
rect 36594 35758 36596 35810
rect 35756 34962 35812 34972
rect 35980 35586 36036 35598
rect 35980 35534 35982 35586
rect 36034 35534 36036 35586
rect 35756 34692 35812 34702
rect 35980 34692 36036 35534
rect 36540 35028 36596 35758
rect 36652 35700 36708 38108
rect 36988 38050 37044 38612
rect 36988 37998 36990 38050
rect 37042 37998 37044 38050
rect 36988 37986 37044 37998
rect 37324 38052 37380 38062
rect 37436 38052 37492 42478
rect 38332 42082 38388 42924
rect 38668 42980 38724 42990
rect 38668 42886 38724 42924
rect 38444 42754 38500 42766
rect 38444 42702 38446 42754
rect 38498 42702 38500 42754
rect 38444 42196 38500 42702
rect 38780 42756 38836 43486
rect 38780 42690 38836 42700
rect 39116 43538 39172 43550
rect 39116 43486 39118 43538
rect 39170 43486 39172 43538
rect 39004 42644 39060 42654
rect 39004 42550 39060 42588
rect 38444 42102 38500 42140
rect 38332 42030 38334 42082
rect 38386 42030 38388 42082
rect 38332 42018 38388 42030
rect 38668 41970 38724 41982
rect 38668 41918 38670 41970
rect 38722 41918 38724 41970
rect 37324 38050 37492 38052
rect 37324 37998 37326 38050
rect 37378 37998 37492 38050
rect 37324 37996 37492 37998
rect 37548 41074 37604 41086
rect 37548 41022 37550 41074
rect 37602 41022 37604 41074
rect 37548 38052 37604 41022
rect 38668 40628 38724 41918
rect 38892 40628 38948 40638
rect 38668 40572 38892 40628
rect 38892 40534 38948 40572
rect 38108 40516 38164 40526
rect 38108 40404 38164 40460
rect 37772 40402 38164 40404
rect 37772 40350 38110 40402
rect 38162 40350 38164 40402
rect 37772 40348 38164 40350
rect 37772 38834 37828 40348
rect 38108 40338 38164 40348
rect 38556 40514 38612 40526
rect 38556 40462 38558 40514
rect 38610 40462 38612 40514
rect 37772 38782 37774 38834
rect 37826 38782 37828 38834
rect 37772 38770 37828 38782
rect 38332 40292 38388 40302
rect 37324 37986 37380 37996
rect 37548 37958 37604 37996
rect 37100 37940 37156 37950
rect 37100 37846 37156 37884
rect 37996 37826 38052 37838
rect 37996 37774 37998 37826
rect 38050 37774 38052 37826
rect 37548 37268 37604 37278
rect 37996 37268 38052 37774
rect 37548 37266 38052 37268
rect 37548 37214 37550 37266
rect 37602 37214 38052 37266
rect 37548 37212 38052 37214
rect 37100 37156 37156 37166
rect 37100 37062 37156 37100
rect 37548 37156 37604 37212
rect 37548 37090 37604 37100
rect 38220 37154 38276 37166
rect 38220 37102 38222 37154
rect 38274 37102 38276 37154
rect 38220 36596 38276 37102
rect 38220 36530 38276 36540
rect 37324 36372 37380 36382
rect 37212 36258 37268 36270
rect 37212 36206 37214 36258
rect 37266 36206 37268 36258
rect 36876 35700 36932 35710
rect 36652 35698 36932 35700
rect 36652 35646 36878 35698
rect 36930 35646 36932 35698
rect 36652 35644 36932 35646
rect 36876 35634 36932 35644
rect 36540 34962 36596 34972
rect 36204 34916 36260 34926
rect 36204 34822 36260 34860
rect 35756 34690 35980 34692
rect 35756 34638 35758 34690
rect 35810 34638 35980 34690
rect 35756 34636 35980 34638
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35756 33236 35812 34636
rect 35980 34598 36036 34636
rect 37100 34692 37156 34702
rect 37100 34598 37156 34636
rect 36988 34468 37044 34478
rect 37212 34468 37268 36206
rect 37324 35698 37380 36316
rect 38332 36036 38388 40236
rect 38444 39732 38500 39742
rect 38444 39638 38500 39676
rect 38556 39284 38612 40462
rect 38556 38724 38612 39228
rect 38556 38668 38724 38724
rect 38668 38612 38948 38668
rect 38892 37940 38948 38612
rect 38892 37938 39060 37940
rect 38892 37886 38894 37938
rect 38946 37886 39060 37938
rect 38892 37884 39060 37886
rect 38892 37874 38948 37884
rect 38556 37828 38612 37838
rect 38556 37826 38724 37828
rect 38556 37774 38558 37826
rect 38610 37774 38724 37826
rect 38556 37772 38724 37774
rect 38556 37762 38612 37772
rect 38668 36482 38724 37772
rect 38668 36430 38670 36482
rect 38722 36430 38724 36482
rect 38668 36418 38724 36430
rect 38780 37826 38836 37838
rect 38780 37774 38782 37826
rect 38834 37774 38836 37826
rect 38780 37156 38836 37774
rect 38780 36372 38836 37100
rect 39004 36708 39060 37884
rect 39004 36642 39060 36652
rect 38892 36596 38948 36606
rect 38892 36502 38948 36540
rect 39116 36482 39172 43486
rect 39340 42756 39396 42766
rect 39340 42642 39396 42700
rect 39340 42590 39342 42642
rect 39394 42590 39396 42642
rect 39340 42578 39396 42590
rect 39116 36430 39118 36482
rect 39170 36430 39172 36482
rect 39116 36418 39172 36430
rect 39228 39396 39284 39406
rect 38780 36316 39060 36372
rect 38332 35980 38612 36036
rect 38444 35810 38500 35822
rect 38444 35758 38446 35810
rect 38498 35758 38500 35810
rect 37324 35646 37326 35698
rect 37378 35646 37380 35698
rect 37324 35634 37380 35646
rect 37884 35698 37940 35710
rect 37884 35646 37886 35698
rect 37938 35646 37940 35698
rect 37884 34914 37940 35646
rect 38220 35700 38276 35710
rect 38220 35606 38276 35644
rect 37884 34862 37886 34914
rect 37938 34862 37940 34914
rect 37044 34412 37268 34468
rect 37324 34802 37380 34814
rect 37324 34750 37326 34802
rect 37378 34750 37380 34802
rect 36652 34018 36708 34030
rect 36652 33966 36654 34018
rect 36706 33966 36708 34018
rect 35756 33170 35812 33180
rect 35868 33908 35924 33918
rect 35308 32564 35364 32574
rect 35308 32470 35364 32508
rect 35532 32340 35588 32350
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35084 31892 35140 31902
rect 34860 27906 34916 27916
rect 34972 30884 35028 30894
rect 34748 27860 34804 27870
rect 34636 27804 34748 27860
rect 33964 27468 34132 27524
rect 33964 27186 34020 27198
rect 33964 27134 33966 27186
rect 34018 27134 34020 27186
rect 33740 27076 33796 27086
rect 33516 26292 33572 26302
rect 33516 24948 33572 26236
rect 33292 24946 33460 24948
rect 33292 24894 33294 24946
rect 33346 24894 33460 24946
rect 33292 24892 33460 24894
rect 33292 24882 33348 24892
rect 32284 24742 32340 24780
rect 32172 24658 32228 24668
rect 33180 24722 33236 24734
rect 33180 24670 33182 24722
rect 33234 24670 33236 24722
rect 32172 24500 32228 24510
rect 32172 24406 32228 24444
rect 33180 23940 33236 24670
rect 33292 24500 33348 24510
rect 33292 24406 33348 24444
rect 32844 23884 33236 23940
rect 33404 24052 33460 24892
rect 33516 24882 33572 24892
rect 33628 25620 33684 25630
rect 31500 19182 31502 19234
rect 31554 19182 31556 19234
rect 31500 19170 31556 19182
rect 31612 19236 31668 19246
rect 32060 19236 32116 20748
rect 32172 23716 32228 23726
rect 32844 23716 32900 23884
rect 33404 23828 33460 23996
rect 32172 23714 32900 23716
rect 32172 23662 32174 23714
rect 32226 23662 32900 23714
rect 32172 23660 32900 23662
rect 32956 23772 33460 23828
rect 32956 23714 33012 23772
rect 32956 23662 32958 23714
rect 33010 23662 33012 23714
rect 32172 20188 32228 23660
rect 32956 23650 33012 23662
rect 33628 23604 33684 25564
rect 33628 23538 33684 23548
rect 33180 21700 33236 21710
rect 33180 21586 33236 21644
rect 33180 21534 33182 21586
rect 33234 21534 33236 21586
rect 33180 21522 33236 21534
rect 33516 21586 33572 21598
rect 33516 21534 33518 21586
rect 33570 21534 33572 21586
rect 33404 21476 33460 21486
rect 33404 21382 33460 21420
rect 33516 20188 33572 21534
rect 33740 20916 33796 27020
rect 33964 26740 34020 27134
rect 33964 26674 34020 26684
rect 34076 26964 34132 27468
rect 34636 27074 34692 27804
rect 34748 27766 34804 27804
rect 34636 27022 34638 27074
rect 34690 27022 34692 27074
rect 34636 27010 34692 27022
rect 34748 27524 34804 27534
rect 33852 26628 33908 26638
rect 33852 24724 33908 26572
rect 33852 24630 33908 24668
rect 33964 23828 34020 23838
rect 34076 23828 34132 26908
rect 34748 26962 34804 27468
rect 34748 26910 34750 26962
rect 34802 26910 34804 26962
rect 34748 26852 34804 26910
rect 34412 26796 34804 26852
rect 34412 26514 34468 26796
rect 34412 26462 34414 26514
rect 34466 26462 34468 26514
rect 34412 26450 34468 26462
rect 34748 26628 34804 26638
rect 34748 26514 34804 26572
rect 34748 26462 34750 26514
rect 34802 26462 34804 26514
rect 34748 26450 34804 26462
rect 34972 26292 35028 30828
rect 35084 30436 35140 31836
rect 35196 31556 35252 31566
rect 35196 31462 35252 31500
rect 35196 30884 35252 30894
rect 35196 30790 35252 30828
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35532 30436 35588 32284
rect 35756 31220 35812 31230
rect 35868 31220 35924 33852
rect 36652 33684 36708 33966
rect 36988 33684 37044 34412
rect 36652 33628 37044 33684
rect 35980 32452 36036 32462
rect 35980 32358 36036 32396
rect 36652 31220 36708 31230
rect 35756 31218 36708 31220
rect 35756 31166 35758 31218
rect 35810 31166 36654 31218
rect 36706 31166 36708 31218
rect 35756 31164 36708 31166
rect 35756 31154 35812 31164
rect 36652 31154 36708 31164
rect 36988 31220 37044 33628
rect 37324 34244 37380 34750
rect 37884 34468 37940 34862
rect 38332 34916 38388 34926
rect 38332 34822 38388 34860
rect 37884 34402 37940 34412
rect 38444 34244 38500 35758
rect 37324 34188 38500 34244
rect 37100 31780 37156 31790
rect 37100 31332 37156 31724
rect 37100 31266 37156 31276
rect 36988 31154 37044 31164
rect 36204 30994 36260 31006
rect 36204 30942 36206 30994
rect 36258 30942 36260 30994
rect 36204 30884 36260 30942
rect 36204 30818 36260 30828
rect 36428 30994 36484 31006
rect 36428 30942 36430 30994
rect 36482 30942 36484 30994
rect 35084 30380 35364 30436
rect 35084 30210 35140 30222
rect 35084 30158 35086 30210
rect 35138 30158 35140 30210
rect 35084 29988 35140 30158
rect 35084 29922 35140 29932
rect 35308 30098 35364 30380
rect 35532 30370 35588 30380
rect 35532 30212 35588 30222
rect 36428 30212 36484 30942
rect 36876 30996 36932 31006
rect 37324 30996 37380 34188
rect 38444 34130 38500 34188
rect 38444 34078 38446 34130
rect 38498 34078 38500 34130
rect 38444 34066 38500 34078
rect 38556 34356 38612 35980
rect 38892 35924 38948 35934
rect 38892 35830 38948 35868
rect 38668 34356 38724 34366
rect 38556 34354 38724 34356
rect 38556 34302 38670 34354
rect 38722 34302 38724 34354
rect 38556 34300 38724 34302
rect 38108 34018 38164 34030
rect 38108 33966 38110 34018
rect 38162 33966 38164 34018
rect 38108 33908 38164 33966
rect 38556 33908 38612 34300
rect 38668 34290 38724 34300
rect 38892 34132 38948 34142
rect 38892 34038 38948 34076
rect 39004 34130 39060 36316
rect 39116 34916 39172 34926
rect 39228 34916 39284 39340
rect 39340 36370 39396 36382
rect 39340 36318 39342 36370
rect 39394 36318 39396 36370
rect 39340 36260 39396 36318
rect 39340 36036 39396 36204
rect 39340 35970 39396 35980
rect 39116 34914 39284 34916
rect 39116 34862 39118 34914
rect 39170 34862 39284 34914
rect 39116 34860 39284 34862
rect 39340 35028 39396 35038
rect 39116 34850 39172 34860
rect 39340 34802 39396 34972
rect 39340 34750 39342 34802
rect 39394 34750 39396 34802
rect 39340 34738 39396 34750
rect 39004 34078 39006 34130
rect 39058 34078 39060 34130
rect 39004 34066 39060 34078
rect 39452 34690 39508 34702
rect 39452 34638 39454 34690
rect 39506 34638 39508 34690
rect 38108 33852 38612 33908
rect 38780 34018 38836 34030
rect 38780 33966 38782 34018
rect 38834 33966 38836 34018
rect 38108 32450 38164 33852
rect 38780 32788 38836 33966
rect 39452 33348 39508 34638
rect 39452 33282 39508 33292
rect 38780 32732 39172 32788
rect 38780 32564 38836 32574
rect 38780 32470 38836 32508
rect 38108 32398 38110 32450
rect 38162 32398 38164 32450
rect 36876 30994 37380 30996
rect 36876 30942 36878 30994
rect 36930 30942 37380 30994
rect 36876 30940 37380 30942
rect 37436 32228 37492 32238
rect 36540 30884 36596 30894
rect 36540 30790 36596 30828
rect 36876 30324 36932 30940
rect 36988 30324 37044 30334
rect 36876 30322 37044 30324
rect 36876 30270 36990 30322
rect 37042 30270 37044 30322
rect 36876 30268 37044 30270
rect 36988 30258 37044 30268
rect 36428 30156 36596 30212
rect 35532 30118 35588 30156
rect 35308 30046 35310 30098
rect 35362 30046 35364 30098
rect 35308 29204 35364 30046
rect 35868 30098 35924 30110
rect 35868 30046 35870 30098
rect 35922 30046 35924 30098
rect 35756 29986 35812 29998
rect 35756 29934 35758 29986
rect 35810 29934 35812 29986
rect 35756 29876 35812 29934
rect 35756 29810 35812 29820
rect 35868 29204 35924 30046
rect 36428 29986 36484 29998
rect 36428 29934 36430 29986
rect 36482 29934 36484 29986
rect 36428 29876 36484 29934
rect 36316 29428 36372 29438
rect 35308 29148 35588 29204
rect 35868 29148 36260 29204
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27860 35252 27870
rect 35084 27804 35196 27860
rect 35084 26908 35140 27804
rect 35196 27794 35252 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 35308 27188 35364 27198
rect 35532 27188 35588 29148
rect 35756 28756 35812 28766
rect 36204 28756 36260 29148
rect 35756 28754 36148 28756
rect 35756 28702 35758 28754
rect 35810 28702 36148 28754
rect 35756 28700 36148 28702
rect 35756 28690 35812 28700
rect 35308 27094 35364 27132
rect 35420 27132 35588 27188
rect 35644 28082 35700 28094
rect 35644 28030 35646 28082
rect 35698 28030 35700 28082
rect 35084 26852 35252 26908
rect 35196 26628 35252 26852
rect 35196 26562 35252 26572
rect 35308 26740 35364 26750
rect 35308 26514 35364 26684
rect 35308 26462 35310 26514
rect 35362 26462 35364 26514
rect 35308 26450 35364 26462
rect 34748 26236 35028 26292
rect 34524 24612 34580 24622
rect 34300 24610 34580 24612
rect 34300 24558 34526 24610
rect 34578 24558 34580 24610
rect 34300 24556 34580 24558
rect 34188 24500 34244 24510
rect 34188 23938 34244 24444
rect 34300 24162 34356 24556
rect 34524 24546 34580 24556
rect 34300 24110 34302 24162
rect 34354 24110 34356 24162
rect 34300 24098 34356 24110
rect 34188 23886 34190 23938
rect 34242 23886 34244 23938
rect 34188 23874 34244 23886
rect 33964 23826 34132 23828
rect 33964 23774 33966 23826
rect 34018 23774 34132 23826
rect 33964 23772 34132 23774
rect 34412 23828 34468 23838
rect 34636 23828 34692 23838
rect 34412 23826 34692 23828
rect 34412 23774 34414 23826
rect 34466 23774 34638 23826
rect 34690 23774 34692 23826
rect 34412 23772 34692 23774
rect 33964 23762 34020 23772
rect 34412 23762 34468 23772
rect 34636 23762 34692 23772
rect 34636 23604 34692 23614
rect 34636 23268 34692 23548
rect 34748 23492 34804 26236
rect 35420 26068 35476 27132
rect 35644 26852 35700 28030
rect 35756 27858 35812 27870
rect 35756 27806 35758 27858
rect 35810 27806 35812 27858
rect 35756 27412 35812 27806
rect 36092 27860 36148 28700
rect 36204 28642 36260 28700
rect 36204 28590 36206 28642
rect 36258 28590 36260 28642
rect 36204 28578 36260 28590
rect 36092 27766 36148 27804
rect 36316 27858 36372 29372
rect 36428 28532 36484 29820
rect 36428 28466 36484 28476
rect 36428 28084 36484 28094
rect 36428 27990 36484 28028
rect 36540 28082 36596 30156
rect 36988 29764 37044 29774
rect 36540 28030 36542 28082
rect 36594 28030 36596 28082
rect 36316 27806 36318 27858
rect 36370 27806 36372 27858
rect 36316 27748 36372 27806
rect 36316 27682 36372 27692
rect 35756 27356 36260 27412
rect 35756 27076 35812 27086
rect 35756 26982 35812 27020
rect 36092 26964 36148 26974
rect 35868 26852 35924 26862
rect 35644 26850 35924 26852
rect 35644 26798 35870 26850
rect 35922 26798 35924 26850
rect 35644 26796 35924 26798
rect 35756 26628 35812 26638
rect 35756 26290 35812 26572
rect 35756 26238 35758 26290
rect 35810 26238 35812 26290
rect 35756 26226 35812 26238
rect 35868 26292 35924 26796
rect 35980 26740 36036 26750
rect 35980 26514 36036 26684
rect 35980 26462 35982 26514
rect 36034 26462 36036 26514
rect 35980 26450 36036 26462
rect 36092 26514 36148 26908
rect 36204 26908 36260 27356
rect 36204 26852 36484 26908
rect 36092 26462 36094 26514
rect 36146 26462 36148 26514
rect 36092 26450 36148 26462
rect 36204 26292 36260 26302
rect 35868 26290 36260 26292
rect 35868 26238 36206 26290
rect 36258 26238 36260 26290
rect 35868 26236 36260 26238
rect 35420 26012 35588 26068
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 35420 25508 35476 25518
rect 35420 25414 35476 25452
rect 34860 24500 34916 24510
rect 34860 23826 34916 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 35196 24164 35252 24174
rect 34860 23774 34862 23826
rect 34914 23774 34916 23826
rect 34860 23762 34916 23774
rect 34972 23826 35028 23838
rect 34972 23774 34974 23826
rect 35026 23774 35028 23826
rect 34972 23716 35028 23774
rect 35028 23660 35140 23716
rect 34972 23650 35028 23660
rect 34748 23436 35028 23492
rect 34748 23268 34804 23278
rect 34188 23266 34804 23268
rect 34188 23214 34750 23266
rect 34802 23214 34804 23266
rect 34188 23212 34804 23214
rect 33964 22372 34020 22382
rect 33964 21924 34020 22316
rect 34188 22370 34244 23212
rect 34748 23202 34804 23212
rect 34748 22930 34804 22942
rect 34748 22878 34750 22930
rect 34802 22878 34804 22930
rect 34188 22318 34190 22370
rect 34242 22318 34244 22370
rect 34188 22306 34244 22318
rect 34636 22372 34692 22382
rect 34748 22372 34804 22878
rect 34636 22370 34804 22372
rect 34636 22318 34638 22370
rect 34690 22318 34804 22370
rect 34636 22316 34804 22318
rect 34636 22306 34692 22316
rect 33964 21858 34020 21868
rect 34076 22146 34132 22158
rect 34076 22094 34078 22146
rect 34130 22094 34132 22146
rect 33852 21700 33908 21710
rect 34076 21700 34132 22094
rect 34860 22148 34916 22158
rect 34860 21810 34916 22092
rect 34860 21758 34862 21810
rect 34914 21758 34916 21810
rect 34860 21746 34916 21758
rect 33852 21698 34132 21700
rect 33852 21646 33854 21698
rect 33906 21646 34132 21698
rect 33852 21644 34132 21646
rect 33852 21634 33908 21644
rect 33852 20916 33908 20926
rect 33740 20914 33908 20916
rect 33740 20862 33854 20914
rect 33906 20862 33908 20914
rect 33740 20860 33908 20862
rect 33852 20188 33908 20860
rect 34972 20188 35028 23436
rect 35084 22370 35140 23660
rect 35196 23378 35252 24108
rect 35196 23326 35198 23378
rect 35250 23326 35252 23378
rect 35196 22930 35252 23326
rect 35196 22878 35198 22930
rect 35250 22878 35252 22930
rect 35196 22866 35252 22878
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 35084 22318 35086 22370
rect 35138 22318 35140 22370
rect 35084 22306 35140 22318
rect 35420 22260 35476 22270
rect 35420 22166 35476 22204
rect 35532 22260 35588 26012
rect 36204 25620 36260 26236
rect 36204 25554 36260 25564
rect 36316 26290 36372 26302
rect 36316 26238 36318 26290
rect 36370 26238 36372 26290
rect 36316 25508 36372 26238
rect 36316 25442 36372 25452
rect 36428 23044 36484 26852
rect 36540 26852 36596 28030
rect 36652 28644 36708 28654
rect 36652 27188 36708 28588
rect 36652 27122 36708 27132
rect 36764 27860 36820 27870
rect 36540 26786 36596 26796
rect 36652 24610 36708 24622
rect 36652 24558 36654 24610
rect 36706 24558 36708 24610
rect 36652 24500 36708 24558
rect 36652 24434 36708 24444
rect 36428 22978 36484 22988
rect 36652 23156 36708 23166
rect 35868 22484 35924 22494
rect 35868 22482 36036 22484
rect 35868 22430 35870 22482
rect 35922 22430 36036 22482
rect 35868 22428 36036 22430
rect 35868 22418 35924 22428
rect 35532 22258 35812 22260
rect 35532 22206 35534 22258
rect 35586 22206 35812 22258
rect 35532 22204 35812 22206
rect 35532 22194 35588 22204
rect 35308 22148 35364 22158
rect 35308 22054 35364 22092
rect 35308 21812 35364 21822
rect 35308 21586 35364 21756
rect 35308 21534 35310 21586
rect 35362 21534 35364 21586
rect 35308 21522 35364 21534
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 32172 20132 32564 20188
rect 33516 20132 33796 20188
rect 33852 20132 34244 20188
rect 32508 19348 32564 20132
rect 32172 19236 32228 19246
rect 32060 19180 32172 19236
rect 31612 19122 31668 19180
rect 32172 19142 32228 19180
rect 32508 19234 32564 19292
rect 32508 19182 32510 19234
rect 32562 19182 32564 19234
rect 32508 19170 32564 19182
rect 33292 19236 33348 19246
rect 33292 19142 33348 19180
rect 31612 19070 31614 19122
rect 31666 19070 31668 19122
rect 31612 19058 31668 19070
rect 31836 19124 31892 19134
rect 31836 19030 31892 19068
rect 32844 19124 32900 19134
rect 32844 19030 32900 19068
rect 32620 19012 32676 19022
rect 32620 18918 32676 18956
rect 32732 19010 32788 19022
rect 32732 18958 32734 19010
rect 32786 18958 32788 19010
rect 31276 18834 31332 18844
rect 32732 17444 32788 18958
rect 33180 18338 33236 18350
rect 33180 18286 33182 18338
rect 33234 18286 33236 18338
rect 32732 17378 32788 17388
rect 32956 17556 33012 17566
rect 33180 17556 33236 18286
rect 33740 18228 33796 20132
rect 33964 19012 34020 19022
rect 33964 18918 34020 18956
rect 33740 18172 34132 18228
rect 33012 17500 33236 17556
rect 33404 17556 33460 17566
rect 32956 17442 33012 17500
rect 33404 17462 33460 17500
rect 32956 17390 32958 17442
rect 33010 17390 33012 17442
rect 32956 17378 33012 17390
rect 33516 17444 33572 17454
rect 32956 17108 33012 17118
rect 32844 16996 32900 17006
rect 32844 16100 32900 16940
rect 32620 16098 32900 16100
rect 32620 16046 32846 16098
rect 32898 16046 32900 16098
rect 32620 16044 32900 16046
rect 31388 15540 31444 15550
rect 31388 15446 31444 15484
rect 32396 15540 32452 15550
rect 32396 15446 32452 15484
rect 31612 15314 31668 15326
rect 31612 15262 31614 15314
rect 31666 15262 31668 15314
rect 31612 15092 31668 15262
rect 31836 15314 31892 15326
rect 31836 15262 31838 15314
rect 31890 15262 31892 15314
rect 31612 15026 31668 15036
rect 31724 15202 31780 15214
rect 31724 15150 31726 15202
rect 31778 15150 31780 15202
rect 31500 14756 31556 14766
rect 31724 14756 31780 15150
rect 31500 14754 31780 14756
rect 31500 14702 31502 14754
rect 31554 14702 31780 14754
rect 31500 14700 31780 14702
rect 31500 14690 31556 14700
rect 31276 14420 31332 14430
rect 31276 14326 31332 14364
rect 31388 14308 31444 14318
rect 31388 14214 31444 14252
rect 31164 13794 31220 13804
rect 31836 13860 31892 15262
rect 32172 15092 32228 15102
rect 31836 13766 31892 13804
rect 31948 14530 32004 14542
rect 31948 14478 31950 14530
rect 32002 14478 32004 14530
rect 31948 13748 32004 14478
rect 32172 14530 32228 15036
rect 32172 14478 32174 14530
rect 32226 14478 32228 14530
rect 32172 14308 32228 14478
rect 32508 14756 32564 14766
rect 32508 14530 32564 14700
rect 32508 14478 32510 14530
rect 32562 14478 32564 14530
rect 32508 14466 32564 14478
rect 32284 14420 32340 14430
rect 32284 14326 32340 14364
rect 32172 13972 32228 14252
rect 32396 14306 32452 14318
rect 32396 14254 32398 14306
rect 32450 14254 32452 14306
rect 32396 14196 32452 14254
rect 32284 13972 32340 13982
rect 32172 13970 32340 13972
rect 32172 13918 32286 13970
rect 32338 13918 32340 13970
rect 32172 13916 32340 13918
rect 32284 13906 32340 13916
rect 31948 13682 32004 13692
rect 32060 13748 32116 13758
rect 32396 13748 32452 14140
rect 32508 13972 32564 13982
rect 32508 13858 32564 13916
rect 32508 13806 32510 13858
rect 32562 13806 32564 13858
rect 32508 13794 32564 13806
rect 32060 13746 32452 13748
rect 32060 13694 32062 13746
rect 32114 13694 32452 13746
rect 32060 13692 32452 13694
rect 32060 13682 32116 13692
rect 31052 13234 31108 13244
rect 31948 13522 32004 13534
rect 32620 13524 32676 16044
rect 32844 16034 32900 16044
rect 32956 16322 33012 17052
rect 33404 16996 33460 17006
rect 33404 16882 33460 16940
rect 33404 16830 33406 16882
rect 33458 16830 33460 16882
rect 33404 16818 33460 16830
rect 33516 16884 33572 17388
rect 33740 16994 33796 18172
rect 34076 17890 34132 18172
rect 34076 17838 34078 17890
rect 34130 17838 34132 17890
rect 34076 17826 34132 17838
rect 33964 17668 34020 17678
rect 34188 17668 34244 20132
rect 34748 20132 35028 20188
rect 34300 19348 34356 19358
rect 34300 19234 34356 19292
rect 34300 19182 34302 19234
rect 34354 19182 34356 19234
rect 34300 19170 34356 19182
rect 34636 19124 34692 19134
rect 34636 19030 34692 19068
rect 34412 19012 34468 19022
rect 34412 18918 34468 18956
rect 33964 17666 34244 17668
rect 33964 17614 33966 17666
rect 34018 17614 34244 17666
rect 33964 17612 34244 17614
rect 33964 17602 34020 17612
rect 33740 16942 33742 16994
rect 33794 16942 33796 16994
rect 33740 16930 33796 16942
rect 34188 16996 34244 17612
rect 34748 17556 34804 20132
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 34860 19348 34916 19358
rect 34860 19234 34916 19292
rect 34860 19182 34862 19234
rect 34914 19182 34916 19234
rect 34860 19170 34916 19182
rect 35308 19236 35364 19246
rect 35756 19236 35812 22204
rect 35980 21698 36036 22428
rect 35980 21646 35982 21698
rect 36034 21646 36036 21698
rect 35980 21634 36036 21646
rect 35364 19180 35812 19236
rect 35196 19124 35252 19134
rect 35196 19030 35252 19068
rect 35308 19122 35364 19180
rect 35308 19070 35310 19122
rect 35362 19070 35364 19122
rect 35308 19058 35364 19070
rect 34972 19010 35028 19022
rect 34972 18958 34974 19010
rect 35026 18958 35028 19010
rect 34972 18452 35028 18958
rect 34972 18386 35028 18396
rect 35084 19010 35140 19022
rect 35084 18958 35086 19010
rect 35138 18958 35140 19010
rect 34748 17490 34804 17500
rect 35084 17444 35140 18958
rect 36428 18564 36484 18574
rect 35420 18450 35476 18462
rect 35420 18398 35422 18450
rect 35474 18398 35476 18450
rect 35420 18340 35476 18398
rect 36092 18452 36148 18462
rect 36092 18358 36148 18396
rect 35420 18274 35476 18284
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 36428 17778 36484 18508
rect 36428 17726 36430 17778
rect 36482 17726 36484 17778
rect 36428 17714 36484 17726
rect 35084 17378 35140 17388
rect 36316 17444 36372 17454
rect 36316 17350 36372 17388
rect 34188 16930 34244 16940
rect 34524 17106 34580 17118
rect 34524 17054 34526 17106
rect 34578 17054 34580 17106
rect 33516 16818 33572 16828
rect 34300 16884 34356 16894
rect 34300 16790 34356 16828
rect 32956 16270 32958 16322
rect 33010 16270 33012 16322
rect 32956 13972 33012 16270
rect 34412 15314 34468 15326
rect 34412 15262 34414 15314
rect 34466 15262 34468 15314
rect 33964 15204 34020 15214
rect 33964 15110 34020 15148
rect 33068 14756 33124 14766
rect 33068 14662 33124 14700
rect 33628 14756 33684 14766
rect 33180 14420 33236 14430
rect 33068 14308 33124 14318
rect 33068 14214 33124 14252
rect 32956 13906 33012 13916
rect 33180 13860 33236 14364
rect 33180 13794 33236 13804
rect 33628 13858 33684 14700
rect 34412 14532 34468 15262
rect 34524 15316 34580 17054
rect 34748 17106 34804 17118
rect 34748 17054 34750 17106
rect 34802 17054 34804 17106
rect 34748 16324 34804 17054
rect 35308 17108 35364 17118
rect 35308 16882 35364 17052
rect 36316 17106 36372 17118
rect 36316 17054 36318 17106
rect 36370 17054 36372 17106
rect 35420 16996 35476 17006
rect 35420 16902 35476 16940
rect 35308 16830 35310 16882
rect 35362 16830 35364 16882
rect 35308 16818 35364 16830
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 34748 16258 34804 16268
rect 36316 16100 36372 17054
rect 36540 17106 36596 17118
rect 36540 17054 36542 17106
rect 36594 17054 36596 17106
rect 36316 16034 36372 16044
rect 36428 16882 36484 16894
rect 36428 16830 36430 16882
rect 36482 16830 36484 16882
rect 36428 16772 36484 16830
rect 34524 15250 34580 15260
rect 34860 15988 34916 15998
rect 34636 15204 34692 15214
rect 34636 15110 34692 15148
rect 34748 14644 34804 14654
rect 34860 14644 34916 15932
rect 36204 15988 36260 15998
rect 35644 15876 35700 15886
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 35644 14756 35700 15820
rect 36204 15876 36260 15932
rect 36428 15876 36484 16716
rect 36204 15820 36484 15876
rect 36204 15314 36260 15820
rect 36204 15262 36206 15314
rect 36258 15262 36260 15314
rect 36204 15250 36260 15262
rect 36540 15314 36596 17054
rect 36540 15262 36542 15314
rect 36594 15262 36596 15314
rect 36540 15204 36596 15262
rect 36540 15138 36596 15148
rect 35644 14754 35812 14756
rect 35644 14702 35646 14754
rect 35698 14702 35812 14754
rect 35644 14700 35812 14702
rect 35644 14690 35700 14700
rect 34748 14642 34916 14644
rect 34748 14590 34750 14642
rect 34802 14590 34916 14642
rect 34748 14588 34916 14590
rect 34748 14578 34804 14588
rect 34412 14466 34468 14476
rect 35308 14420 35364 14430
rect 35308 14326 35364 14364
rect 33852 13972 33908 13982
rect 33852 13878 33908 13916
rect 33628 13806 33630 13858
rect 33682 13806 33684 13858
rect 33628 13794 33684 13806
rect 35532 13746 35588 13758
rect 35532 13694 35534 13746
rect 35586 13694 35588 13746
rect 31948 13470 31950 13522
rect 32002 13470 32004 13522
rect 28588 12982 28644 13020
rect 27692 12350 27694 12402
rect 27746 12350 27748 12402
rect 27692 12338 27748 12350
rect 28812 12404 28868 12414
rect 28812 12310 28868 12348
rect 29260 12404 29316 12414
rect 27580 12238 27582 12290
rect 27634 12238 27636 12290
rect 27580 12226 27636 12238
rect 27244 10722 27300 12124
rect 27356 12178 27412 12190
rect 27356 12126 27358 12178
rect 27410 12126 27412 12178
rect 27356 11956 27412 12126
rect 29260 12178 29316 12348
rect 29260 12126 29262 12178
rect 29314 12126 29316 12178
rect 29260 12114 29316 12126
rect 29932 12066 29988 12078
rect 29932 12014 29934 12066
rect 29986 12014 29988 12066
rect 27692 11956 27748 11966
rect 27356 11954 27748 11956
rect 27356 11902 27694 11954
rect 27746 11902 27748 11954
rect 27356 11900 27748 11902
rect 27692 11890 27748 11900
rect 29932 11508 29988 12014
rect 31948 11788 32004 13470
rect 32060 13468 32676 13524
rect 33964 13522 34020 13534
rect 33964 13470 33966 13522
rect 34018 13470 34020 13522
rect 32060 12068 32116 13468
rect 33068 12740 33124 12750
rect 32060 12066 32452 12068
rect 32060 12014 32062 12066
rect 32114 12014 32452 12066
rect 32060 12012 32452 12014
rect 32060 12002 32116 12012
rect 29932 11442 29988 11452
rect 31724 11732 32004 11788
rect 31500 11394 31556 11406
rect 31500 11342 31502 11394
rect 31554 11342 31556 11394
rect 28028 11284 28084 11294
rect 27356 10948 27412 10958
rect 27356 10834 27412 10892
rect 27356 10782 27358 10834
rect 27410 10782 27412 10834
rect 27356 10770 27412 10782
rect 27916 10948 27972 10958
rect 27916 10834 27972 10892
rect 27916 10782 27918 10834
rect 27970 10782 27972 10834
rect 27916 10770 27972 10782
rect 27244 10670 27246 10722
rect 27298 10670 27300 10722
rect 27244 10658 27300 10670
rect 27356 10386 27412 10398
rect 27356 10334 27358 10386
rect 27410 10334 27412 10386
rect 27356 9826 27412 10334
rect 27356 9774 27358 9826
rect 27410 9774 27412 9826
rect 27356 9762 27412 9774
rect 28028 9826 28084 11228
rect 31500 11284 31556 11342
rect 31724 11394 31780 11732
rect 31836 11508 31892 11518
rect 31836 11414 31892 11452
rect 31724 11342 31726 11394
rect 31778 11342 31780 11394
rect 31724 11330 31780 11342
rect 31500 11218 31556 11228
rect 31948 11284 32004 11294
rect 32172 11284 32228 11294
rect 31948 11282 32228 11284
rect 31948 11230 31950 11282
rect 32002 11230 32174 11282
rect 32226 11230 32228 11282
rect 31948 11228 32228 11230
rect 31948 11218 32004 11228
rect 32172 11218 32228 11228
rect 32396 11282 32452 12012
rect 33068 12066 33124 12684
rect 33068 12014 33070 12066
rect 33122 12014 33124 12066
rect 33068 12002 33124 12014
rect 33964 11956 34020 13470
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35532 12740 35588 13694
rect 35756 13634 35812 14700
rect 35756 13582 35758 13634
rect 35810 13582 35812 13634
rect 35756 13570 35812 13582
rect 35868 14532 35924 14542
rect 35644 13188 35700 13198
rect 35644 12962 35700 13132
rect 35644 12910 35646 12962
rect 35698 12910 35700 12962
rect 35644 12898 35700 12910
rect 35532 12674 35588 12684
rect 35868 12740 35924 14476
rect 36204 13634 36260 13646
rect 36204 13582 36206 13634
rect 36258 13582 36260 13634
rect 36204 12962 36260 13582
rect 36204 12910 36206 12962
rect 36258 12910 36260 12962
rect 36204 12898 36260 12910
rect 35868 12646 35924 12684
rect 35980 12738 36036 12750
rect 35980 12686 35982 12738
rect 36034 12686 36036 12738
rect 33964 11890 34020 11900
rect 34972 12404 35028 12414
rect 35980 12404 36036 12686
rect 36092 12740 36148 12750
rect 36092 12646 36148 12684
rect 35980 12348 36372 12404
rect 32396 11230 32398 11282
rect 32450 11230 32452 11282
rect 32396 11218 32452 11230
rect 32508 11282 32564 11294
rect 32508 11230 32510 11282
rect 32562 11230 32564 11282
rect 28028 9774 28030 9826
rect 28082 9774 28084 9826
rect 28028 9762 28084 9774
rect 29820 10948 29876 10958
rect 27804 9714 27860 9726
rect 27804 9662 27806 9714
rect 27858 9662 27860 9714
rect 27692 9602 27748 9614
rect 27692 9550 27694 9602
rect 27746 9550 27748 9602
rect 27692 9154 27748 9550
rect 27692 9102 27694 9154
rect 27746 9102 27748 9154
rect 27692 9090 27748 9102
rect 27020 9042 27076 9054
rect 27020 8990 27022 9042
rect 27074 8990 27076 9042
rect 27020 8484 27076 8990
rect 27020 8418 27076 8428
rect 26796 6862 26798 6914
rect 26850 6862 26852 6914
rect 26796 6850 26852 6862
rect 27244 7586 27300 7598
rect 27244 7534 27246 7586
rect 27298 7534 27300 7586
rect 26908 6580 26964 6590
rect 27244 6580 27300 7534
rect 27580 7588 27636 7598
rect 27580 7494 27636 7532
rect 27804 6690 27860 9662
rect 29372 8932 29428 8942
rect 29036 8036 29092 8046
rect 29036 7698 29092 7980
rect 29036 7646 29038 7698
rect 29090 7646 29092 7698
rect 29036 7634 29092 7646
rect 29372 7698 29428 8876
rect 29820 8930 29876 10892
rect 31500 10164 31556 10174
rect 29820 8878 29822 8930
rect 29874 8878 29876 8930
rect 29820 8866 29876 8878
rect 30268 10052 30324 10062
rect 30268 9938 30324 9996
rect 30268 9886 30270 9938
rect 30322 9886 30324 9938
rect 30268 8428 30324 9886
rect 30716 9604 30772 9614
rect 31164 9604 31220 9614
rect 30716 9602 31220 9604
rect 30716 9550 30718 9602
rect 30770 9550 31166 9602
rect 31218 9550 31220 9602
rect 30716 9548 31220 9550
rect 30716 9538 30772 9548
rect 31164 9492 31220 9548
rect 31164 9426 31220 9436
rect 31500 9268 31556 10108
rect 32508 9828 32564 11230
rect 32508 9762 32564 9772
rect 32732 11284 32788 11294
rect 32732 9826 32788 11228
rect 34972 10164 35028 12348
rect 36316 12290 36372 12348
rect 36316 12238 36318 12290
rect 36370 12238 36372 12290
rect 36316 12226 36372 12238
rect 36540 12290 36596 12302
rect 36540 12238 36542 12290
rect 36594 12238 36596 12290
rect 35980 12180 36036 12190
rect 35196 12068 35252 12078
rect 35196 11974 35252 12012
rect 35420 11956 35476 11966
rect 35476 11900 35588 11956
rect 35420 11890 35476 11900
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 34972 10098 35028 10108
rect 34860 10052 34916 10062
rect 34860 9938 34916 9996
rect 34860 9886 34862 9938
rect 34914 9886 34916 9938
rect 34860 9874 34916 9886
rect 35420 10052 35476 10062
rect 35532 10052 35588 11900
rect 35980 11172 36036 12124
rect 36428 12068 36484 12078
rect 36428 11974 36484 12012
rect 36540 11844 36596 12238
rect 36540 11778 36596 11788
rect 36204 11172 36260 11182
rect 35980 11170 36260 11172
rect 35980 11118 36206 11170
rect 36258 11118 36260 11170
rect 35980 11116 36260 11118
rect 35420 10050 35588 10052
rect 35420 9998 35422 10050
rect 35474 9998 35588 10050
rect 35420 9996 35588 9998
rect 35868 10052 35924 10062
rect 32732 9774 32734 9826
rect 32786 9774 32788 9826
rect 32732 9762 32788 9774
rect 33404 9826 33460 9838
rect 33404 9774 33406 9826
rect 33458 9774 33460 9826
rect 32956 9716 33012 9726
rect 32956 9622 33012 9660
rect 30940 9266 31556 9268
rect 30940 9214 31502 9266
rect 31554 9214 31556 9266
rect 30940 9212 31556 9214
rect 30940 9042 30996 9212
rect 31500 9202 31556 9212
rect 33068 9602 33124 9614
rect 33068 9550 33070 9602
rect 33122 9550 33124 9602
rect 30940 8990 30942 9042
rect 30994 8990 30996 9042
rect 30940 8978 30996 8990
rect 30716 8932 30772 8942
rect 30716 8838 30772 8876
rect 30604 8820 30660 8830
rect 30268 8372 30436 8428
rect 30156 8036 30212 8046
rect 30044 8034 30212 8036
rect 30044 7982 30158 8034
rect 30210 7982 30212 8034
rect 30044 7980 30212 7982
rect 29708 7700 29764 7710
rect 29372 7646 29374 7698
rect 29426 7646 29428 7698
rect 27804 6638 27806 6690
rect 27858 6638 27860 6690
rect 27804 6626 27860 6638
rect 29372 6692 29428 7646
rect 29596 7644 29708 7700
rect 29484 6692 29540 6702
rect 29372 6690 29540 6692
rect 29372 6638 29486 6690
rect 29538 6638 29540 6690
rect 29372 6636 29540 6638
rect 29484 6626 29540 6636
rect 27468 6580 27524 6590
rect 26908 6578 27524 6580
rect 26908 6526 26910 6578
rect 26962 6526 27470 6578
rect 27522 6526 27524 6578
rect 26908 6524 27524 6526
rect 26908 6514 26964 6524
rect 26796 6468 26852 6478
rect 26796 6374 26852 6412
rect 27468 6132 27524 6524
rect 27580 6466 27636 6478
rect 27580 6414 27582 6466
rect 27634 6414 27636 6466
rect 27580 6244 27636 6414
rect 29260 6466 29316 6478
rect 29260 6414 29262 6466
rect 29314 6414 29316 6466
rect 27636 6188 27972 6244
rect 27580 6178 27636 6188
rect 27468 6066 27524 6076
rect 27916 5124 27972 6188
rect 28140 5908 28196 5918
rect 27916 5122 28084 5124
rect 27916 5070 27918 5122
rect 27970 5070 28084 5122
rect 27916 5068 28084 5070
rect 27916 5058 27972 5068
rect 26348 4274 26404 4284
rect 28028 4228 28084 5068
rect 28140 5010 28196 5852
rect 29260 5908 29316 6414
rect 29260 5842 29316 5852
rect 29596 5684 29652 7644
rect 29708 7634 29764 7644
rect 30044 7476 30100 7980
rect 30156 7970 30212 7980
rect 30268 7700 30324 7710
rect 30268 7606 30324 7644
rect 30044 7382 30100 7420
rect 29372 5628 29652 5684
rect 29708 5908 29764 5918
rect 29372 5236 29428 5628
rect 28588 5234 29428 5236
rect 28588 5182 29374 5234
rect 29426 5182 29428 5234
rect 28588 5180 29428 5182
rect 28252 5124 28308 5134
rect 28252 5030 28308 5068
rect 28588 5122 28644 5180
rect 29372 5170 29428 5180
rect 29596 5236 29652 5246
rect 29596 5142 29652 5180
rect 28588 5070 28590 5122
rect 28642 5070 28644 5122
rect 28588 5058 28644 5070
rect 29708 5122 29764 5852
rect 29708 5070 29710 5122
rect 29762 5070 29764 5122
rect 29708 5058 29764 5070
rect 30156 5348 30212 5358
rect 30156 5122 30212 5292
rect 30380 5236 30436 8372
rect 30492 8260 30548 8270
rect 30604 8260 30660 8764
rect 30492 8258 30660 8260
rect 30492 8206 30494 8258
rect 30546 8206 30660 8258
rect 30492 8204 30660 8206
rect 31276 8484 31332 8494
rect 33068 8428 33124 9550
rect 33404 8932 33460 9774
rect 33852 9828 33908 9838
rect 33852 9734 33908 9772
rect 35308 9828 35364 9838
rect 33516 9716 33572 9726
rect 34636 9716 34692 9726
rect 33516 9622 33572 9660
rect 34524 9714 34692 9716
rect 34524 9662 34638 9714
rect 34690 9662 34692 9714
rect 34524 9660 34692 9662
rect 33740 9602 33796 9614
rect 33740 9550 33742 9602
rect 33794 9550 33796 9602
rect 33740 9492 33796 9550
rect 34524 9492 34580 9660
rect 34636 9650 34692 9660
rect 35308 9602 35364 9772
rect 35308 9550 35310 9602
rect 35362 9550 35364 9602
rect 35308 9538 35364 9550
rect 33740 9436 34580 9492
rect 33404 8866 33460 8876
rect 31276 8260 31332 8428
rect 32396 8372 33124 8428
rect 32396 8370 32452 8372
rect 32396 8318 32398 8370
rect 32450 8318 32452 8370
rect 32396 8306 32452 8318
rect 34524 8370 34580 9436
rect 35420 9154 35476 9996
rect 35644 9828 35700 9838
rect 35644 9826 35812 9828
rect 35644 9774 35646 9826
rect 35698 9774 35812 9826
rect 35644 9772 35812 9774
rect 35644 9762 35700 9772
rect 35644 9268 35700 9278
rect 35644 9174 35700 9212
rect 35420 9102 35422 9154
rect 35474 9102 35476 9154
rect 35420 9090 35476 9102
rect 35532 8932 35588 8942
rect 35532 8838 35588 8876
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 34524 8318 34526 8370
rect 34578 8318 34580 8370
rect 34524 8306 34580 8318
rect 31612 8260 31668 8270
rect 31276 8258 31668 8260
rect 31276 8206 31278 8258
rect 31330 8206 31614 8258
rect 31666 8206 31668 8258
rect 31276 8204 31668 8206
rect 30492 8194 30548 8204
rect 31276 8194 31332 8204
rect 31612 8194 31668 8204
rect 32284 7700 32340 7710
rect 32172 6804 32228 6814
rect 32172 6710 32228 6748
rect 32284 6690 32340 7644
rect 33180 7700 33236 7710
rect 33180 7606 33236 7644
rect 35756 7476 35812 9772
rect 35868 9266 35924 9996
rect 35980 9716 36036 9726
rect 35980 9622 36036 9660
rect 35868 9214 35870 9266
rect 35922 9214 35924 9266
rect 35868 9202 35924 9214
rect 36092 8428 36148 11116
rect 36204 11106 36260 11116
rect 36204 10388 36260 10398
rect 36204 10050 36260 10332
rect 36204 9998 36206 10050
rect 36258 9998 36260 10050
rect 36204 9986 36260 9998
rect 36652 8428 36708 23100
rect 36764 16772 36820 27804
rect 36988 24164 37044 29708
rect 37436 28084 37492 32172
rect 37548 31556 37604 31566
rect 38108 31556 38164 32398
rect 37548 31554 37716 31556
rect 37548 31502 37550 31554
rect 37602 31502 37716 31554
rect 37548 31500 37716 31502
rect 37548 31490 37604 31500
rect 37548 31332 37604 31342
rect 37548 31106 37604 31276
rect 37548 31054 37550 31106
rect 37602 31054 37604 31106
rect 37548 31042 37604 31054
rect 37660 31108 37716 31500
rect 38108 31490 38164 31500
rect 38892 31666 38948 31678
rect 38892 31614 38894 31666
rect 38946 31614 38948 31666
rect 38668 31220 38724 31230
rect 38444 31218 38724 31220
rect 38444 31166 38670 31218
rect 38722 31166 38724 31218
rect 38444 31164 38724 31166
rect 37772 31108 37828 31118
rect 38444 31108 38500 31164
rect 38668 31154 38724 31164
rect 38892 31218 38948 31614
rect 38892 31166 38894 31218
rect 38946 31166 38948 31218
rect 38892 31154 38948 31166
rect 39004 31554 39060 31566
rect 39004 31502 39006 31554
rect 39058 31502 39060 31554
rect 37660 31052 37772 31108
rect 37772 31014 37828 31052
rect 38220 31052 38500 31108
rect 37884 30996 37940 31006
rect 37884 30902 37940 30940
rect 37996 30994 38052 31006
rect 37996 30942 37998 30994
rect 38050 30942 38052 30994
rect 37996 30100 38052 30942
rect 37996 30034 38052 30044
rect 38108 30994 38164 31006
rect 38108 30942 38110 30994
rect 38162 30942 38164 30994
rect 37548 29988 37604 29998
rect 37548 29986 37716 29988
rect 37548 29934 37550 29986
rect 37602 29934 37716 29986
rect 37548 29932 37716 29934
rect 37548 29922 37604 29932
rect 37548 28868 37604 28878
rect 37548 28642 37604 28812
rect 37660 28756 37716 29932
rect 38108 29876 38164 30942
rect 38220 30324 38276 31052
rect 38556 30996 38612 31006
rect 38220 30210 38276 30268
rect 38220 30158 38222 30210
rect 38274 30158 38276 30210
rect 38220 30146 38276 30158
rect 38332 30994 38612 30996
rect 38332 30942 38558 30994
rect 38610 30942 38612 30994
rect 38332 30940 38612 30942
rect 37660 28690 37716 28700
rect 37772 29820 38164 29876
rect 37548 28590 37550 28642
rect 37602 28590 37604 28642
rect 37548 28578 37604 28590
rect 37772 28642 37828 29820
rect 37884 29652 37940 29662
rect 37884 29558 37940 29596
rect 38220 29540 38276 29550
rect 38332 29540 38388 30940
rect 38556 30930 38612 30940
rect 39004 30324 39060 31502
rect 39116 31220 39172 32732
rect 39228 32562 39284 32574
rect 39228 32510 39230 32562
rect 39282 32510 39284 32562
rect 39228 31778 39284 32510
rect 39452 32452 39508 32462
rect 39452 32358 39508 32396
rect 39228 31726 39230 31778
rect 39282 31726 39284 31778
rect 39228 31714 39284 31726
rect 39228 31220 39284 31230
rect 39116 31218 39284 31220
rect 39116 31166 39230 31218
rect 39282 31166 39284 31218
rect 39116 31164 39284 31166
rect 39228 31154 39284 31164
rect 39116 30996 39172 31006
rect 39116 30902 39172 30940
rect 39228 30772 39284 30782
rect 39228 30678 39284 30716
rect 39004 30258 39060 30268
rect 39452 30100 39508 30110
rect 38220 29538 38388 29540
rect 38220 29486 38222 29538
rect 38274 29486 38388 29538
rect 38220 29484 38388 29486
rect 38444 29652 38500 29662
rect 38444 29538 38500 29596
rect 39004 29652 39060 29662
rect 39452 29652 39508 30044
rect 39564 29764 39620 44044
rect 39676 43988 39732 46508
rect 39788 45890 39844 45902
rect 39788 45838 39790 45890
rect 39842 45838 39844 45890
rect 39788 45668 39844 45838
rect 39788 45602 39844 45612
rect 40012 45108 40068 46620
rect 40236 46674 40292 46686
rect 40236 46622 40238 46674
rect 40290 46622 40292 46674
rect 40236 45892 40292 46622
rect 40236 45826 40292 45836
rect 40572 45892 40628 45902
rect 40572 45778 40628 45836
rect 40572 45726 40574 45778
rect 40626 45726 40628 45778
rect 40572 45714 40628 45726
rect 40236 45668 40292 45678
rect 40236 45574 40292 45612
rect 39676 43932 39844 43988
rect 39676 42644 39732 42654
rect 39676 42550 39732 42588
rect 39788 37044 39844 43932
rect 39900 42644 39956 42654
rect 39900 42082 39956 42588
rect 40012 42194 40068 45052
rect 40012 42142 40014 42194
rect 40066 42142 40068 42194
rect 40012 42130 40068 42142
rect 40348 42756 40404 42766
rect 39900 42030 39902 42082
rect 39954 42030 39956 42082
rect 39900 42018 39956 42030
rect 40236 41970 40292 41982
rect 40236 41918 40238 41970
rect 40290 41918 40292 41970
rect 40236 41076 40292 41918
rect 40236 41010 40292 41020
rect 39788 36978 39844 36988
rect 39900 40572 40180 40628
rect 39900 39732 39956 40572
rect 40124 40514 40180 40572
rect 40124 40462 40126 40514
rect 40178 40462 40180 40514
rect 40124 40450 40180 40462
rect 40012 40404 40068 40414
rect 40012 40310 40068 40348
rect 40236 40404 40292 40414
rect 40124 40180 40180 40190
rect 40236 40180 40292 40348
rect 40124 40178 40292 40180
rect 40124 40126 40126 40178
rect 40178 40126 40292 40178
rect 40124 40124 40292 40126
rect 40124 40114 40180 40124
rect 39676 36708 39732 36718
rect 39676 32674 39732 36652
rect 39788 36260 39844 36270
rect 39788 36166 39844 36204
rect 39788 34356 39844 34366
rect 39900 34356 39956 39676
rect 40348 39620 40404 42700
rect 40796 42420 40852 50876
rect 41244 50708 41300 50718
rect 41132 50706 41300 50708
rect 41132 50654 41246 50706
rect 41298 50654 41300 50706
rect 41132 50652 41300 50654
rect 41132 49252 41188 50652
rect 41244 50642 41300 50652
rect 48300 50708 48356 50718
rect 48300 50706 48468 50708
rect 48300 50654 48302 50706
rect 48354 50654 48468 50706
rect 48300 50652 48468 50654
rect 48300 50642 48356 50652
rect 44156 50594 44212 50606
rect 44156 50542 44158 50594
rect 44210 50542 44212 50594
rect 43372 50484 43428 50494
rect 42140 50482 43428 50484
rect 42140 50430 43374 50482
rect 43426 50430 43428 50482
rect 42140 50428 43428 50430
rect 42028 49922 42084 49934
rect 42028 49870 42030 49922
rect 42082 49870 42084 49922
rect 41804 49588 41860 49598
rect 40908 49028 40964 49038
rect 40908 48934 40964 48972
rect 41132 49026 41188 49196
rect 41244 49586 41860 49588
rect 41244 49534 41806 49586
rect 41858 49534 41860 49586
rect 41244 49532 41860 49534
rect 41244 49138 41300 49532
rect 41804 49522 41860 49532
rect 41244 49086 41246 49138
rect 41298 49086 41300 49138
rect 41244 49074 41300 49086
rect 41132 48974 41134 49026
rect 41186 48974 41188 49026
rect 41132 48962 41188 48974
rect 41356 48916 41412 48926
rect 41356 48822 41412 48860
rect 41580 48916 41636 48926
rect 41580 48914 41748 48916
rect 41580 48862 41582 48914
rect 41634 48862 41748 48914
rect 41580 48860 41748 48862
rect 41580 48850 41636 48860
rect 41020 48132 41076 48142
rect 41020 48038 41076 48076
rect 41580 47460 41636 47470
rect 41580 47366 41636 47404
rect 41692 47236 41748 48860
rect 42028 48468 42084 49870
rect 42140 49698 42196 50428
rect 43372 50418 43428 50428
rect 44156 50484 44212 50542
rect 45500 50594 45556 50606
rect 45500 50542 45502 50594
rect 45554 50542 45556 50594
rect 44156 50418 44212 50428
rect 44940 50484 44996 50494
rect 45500 50484 45556 50542
rect 44996 50428 45556 50484
rect 44940 50390 44996 50428
rect 42140 49646 42142 49698
rect 42194 49646 42196 49698
rect 42140 49634 42196 49646
rect 42140 48468 42196 48478
rect 42028 48466 42868 48468
rect 42028 48414 42142 48466
rect 42194 48414 42868 48466
rect 42028 48412 42868 48414
rect 42140 48402 42196 48412
rect 42476 48242 42532 48254
rect 42476 48190 42478 48242
rect 42530 48190 42532 48242
rect 41804 48132 41860 48142
rect 41804 48038 41860 48076
rect 42476 48132 42532 48190
rect 41916 47348 41972 47358
rect 41916 47254 41972 47292
rect 42252 47346 42308 47358
rect 42252 47294 42254 47346
rect 42306 47294 42308 47346
rect 41804 47236 41860 47246
rect 41692 47180 41804 47236
rect 41804 47142 41860 47180
rect 42028 47234 42084 47246
rect 42028 47182 42030 47234
rect 42082 47182 42084 47234
rect 41132 45892 41188 45902
rect 41132 45330 41188 45836
rect 42028 45892 42084 47182
rect 42252 46452 42308 47294
rect 42476 46676 42532 48076
rect 42700 47348 42756 47358
rect 42700 47254 42756 47292
rect 42812 47348 42868 48412
rect 42924 48242 42980 48254
rect 42924 48190 42926 48242
rect 42978 48190 42980 48242
rect 42924 48132 42980 48190
rect 43596 48132 43652 48142
rect 42924 48066 42980 48076
rect 43036 48130 43652 48132
rect 43036 48078 43598 48130
rect 43650 48078 43652 48130
rect 43036 48076 43652 48078
rect 43036 47682 43092 48076
rect 43596 48066 43652 48076
rect 45500 48132 45556 50428
rect 46172 50484 46228 50494
rect 46172 50482 46900 50484
rect 46172 50430 46174 50482
rect 46226 50430 46900 50482
rect 46172 50428 46900 50430
rect 46172 50418 46228 50428
rect 46732 48914 46788 48926
rect 46732 48862 46734 48914
rect 46786 48862 46788 48914
rect 46396 48804 46452 48814
rect 46396 48710 46452 48748
rect 46508 48242 46564 48254
rect 46508 48190 46510 48242
rect 46562 48190 46564 48242
rect 45500 48066 45556 48076
rect 45724 48130 45780 48142
rect 45724 48078 45726 48130
rect 45778 48078 45780 48130
rect 43036 47630 43038 47682
rect 43090 47630 43092 47682
rect 43036 47618 43092 47630
rect 42924 47348 42980 47358
rect 42812 47346 42980 47348
rect 42812 47294 42926 47346
rect 42978 47294 42980 47346
rect 42812 47292 42980 47294
rect 42476 46610 42532 46620
rect 42252 46386 42308 46396
rect 42812 46116 42868 47292
rect 42924 47282 42980 47292
rect 45724 47236 45780 48078
rect 46172 48132 46228 48142
rect 46172 48038 46228 48076
rect 45724 46676 45780 47180
rect 45500 46620 45780 46676
rect 46172 47236 46228 47246
rect 46508 47236 46564 48190
rect 46732 47348 46788 48862
rect 46844 48466 46900 50428
rect 48300 49700 48356 49710
rect 48188 49644 48300 49700
rect 47068 49138 47124 49150
rect 47068 49086 47070 49138
rect 47122 49086 47124 49138
rect 46956 48804 47012 48814
rect 46956 48710 47012 48748
rect 46844 48414 46846 48466
rect 46898 48414 46900 48466
rect 46844 48402 46900 48414
rect 47068 48354 47124 49086
rect 47180 48916 47236 48926
rect 47180 48822 47236 48860
rect 47068 48302 47070 48354
rect 47122 48302 47124 48354
rect 47068 48290 47124 48302
rect 48188 48804 48244 49644
rect 48300 49606 48356 49644
rect 48412 48916 48468 50652
rect 48748 50372 48804 50382
rect 48748 50278 48804 50316
rect 49644 50034 49700 51324
rect 49980 51378 50036 51390
rect 49980 51326 49982 51378
rect 50034 51326 50036 51378
rect 49644 49982 49646 50034
rect 49698 49982 49700 50034
rect 49644 49970 49700 49982
rect 49756 51268 49812 51278
rect 49980 51268 50036 51326
rect 49756 51266 50036 51268
rect 49756 51214 49758 51266
rect 49810 51214 50036 51266
rect 49756 51212 50036 51214
rect 50428 51378 50484 51390
rect 50428 51326 50430 51378
rect 50482 51326 50484 51378
rect 50428 51268 50484 51326
rect 50652 51380 50708 51390
rect 50652 51286 50708 51324
rect 48748 49812 48804 49822
rect 48748 49810 49140 49812
rect 48748 49758 48750 49810
rect 48802 49758 49140 49810
rect 48748 49756 49140 49758
rect 48748 49746 48804 49756
rect 48972 49586 49028 49598
rect 48972 49534 48974 49586
rect 49026 49534 49028 49586
rect 48748 49028 48804 49038
rect 48748 48934 48804 48972
rect 48972 49026 49028 49534
rect 48972 48974 48974 49026
rect 49026 48974 49028 49026
rect 48972 48916 49028 48974
rect 49084 49028 49140 49756
rect 49196 49700 49252 49710
rect 49196 49606 49252 49644
rect 49756 49252 49812 51212
rect 49980 50372 50036 50382
rect 49980 49700 50036 50316
rect 50428 50036 50484 51212
rect 51100 50818 51156 51548
rect 51212 51380 51268 51390
rect 51212 51286 51268 51324
rect 51436 51378 51492 51390
rect 51436 51326 51438 51378
rect 51490 51326 51492 51378
rect 51100 50766 51102 50818
rect 51154 50766 51156 50818
rect 51100 50754 51156 50766
rect 51324 51266 51380 51278
rect 51324 51214 51326 51266
rect 51378 51214 51380 51266
rect 50556 50204 50820 50214
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50556 50138 50820 50148
rect 50428 49980 50596 50036
rect 50316 49810 50372 49822
rect 50316 49758 50318 49810
rect 50370 49758 50372 49810
rect 50316 49700 50372 49758
rect 49980 49698 50372 49700
rect 49980 49646 49982 49698
rect 50034 49646 50372 49698
rect 49980 49644 50372 49646
rect 49980 49634 50036 49644
rect 49644 49196 49812 49252
rect 49196 49028 49252 49038
rect 49084 49026 49252 49028
rect 49084 48974 49198 49026
rect 49250 48974 49252 49026
rect 49084 48972 49252 48974
rect 48412 48850 48468 48860
rect 48860 48860 48972 48916
rect 46844 48244 46900 48254
rect 46844 48150 46900 48188
rect 46732 47282 46788 47292
rect 47180 48132 47236 48142
rect 46172 47234 46564 47236
rect 46172 47182 46174 47234
rect 46226 47182 46564 47234
rect 46172 47180 46564 47182
rect 44156 46564 44212 46574
rect 42700 46060 42868 46116
rect 42924 46452 42980 46462
rect 42364 46004 42420 46014
rect 42364 46002 42532 46004
rect 42364 45950 42366 46002
rect 42418 45950 42532 46002
rect 42364 45948 42532 45950
rect 42364 45938 42420 45948
rect 42028 45798 42084 45836
rect 41132 45278 41134 45330
rect 41186 45278 41188 45330
rect 41132 45266 41188 45278
rect 41468 45780 41524 45790
rect 40908 45108 40964 45118
rect 40908 45014 40964 45052
rect 41356 45106 41412 45118
rect 41356 45054 41358 45106
rect 41410 45054 41412 45106
rect 41244 44994 41300 45006
rect 41244 44942 41246 44994
rect 41298 44942 41300 44994
rect 41020 42644 41076 42654
rect 41020 42642 41188 42644
rect 41020 42590 41022 42642
rect 41074 42590 41188 42642
rect 41020 42588 41188 42590
rect 41020 42578 41076 42588
rect 40796 42364 41076 42420
rect 40908 41970 40964 41982
rect 40908 41918 40910 41970
rect 40962 41918 40964 41970
rect 40572 40964 40628 40974
rect 40908 40964 40964 41918
rect 41020 41748 41076 42364
rect 41132 42194 41188 42588
rect 41132 42142 41134 42194
rect 41186 42142 41188 42194
rect 41132 42130 41188 42142
rect 41244 41970 41300 44942
rect 41356 44884 41412 45054
rect 41468 45106 41524 45724
rect 41468 45054 41470 45106
rect 41522 45054 41524 45106
rect 41468 45042 41524 45054
rect 41804 45778 41860 45790
rect 41804 45726 41806 45778
rect 41858 45726 41860 45778
rect 41804 44884 41860 45726
rect 42364 45780 42420 45790
rect 42364 45686 42420 45724
rect 42252 45666 42308 45678
rect 42252 45614 42254 45666
rect 42306 45614 42308 45666
rect 42252 45332 42308 45614
rect 42476 45332 42532 45948
rect 42700 45556 42756 46060
rect 42924 45892 42980 46396
rect 44156 46114 44212 46508
rect 44156 46062 44158 46114
rect 44210 46062 44212 46114
rect 44156 46050 44212 46062
rect 44380 46562 44436 46574
rect 44380 46510 44382 46562
rect 44434 46510 44436 46562
rect 44380 46452 44436 46510
rect 43036 45892 43092 45902
rect 42924 45890 43092 45892
rect 42924 45838 43038 45890
rect 43090 45838 43092 45890
rect 42924 45836 43092 45838
rect 43036 45826 43092 45836
rect 43260 45892 43316 45902
rect 43260 45798 43316 45836
rect 43372 45890 43428 45902
rect 43372 45838 43374 45890
rect 43426 45838 43428 45890
rect 43148 45780 43204 45790
rect 43148 45686 43204 45724
rect 42924 45668 42980 45678
rect 42924 45574 42980 45612
rect 42700 45490 42756 45500
rect 43148 45556 43204 45566
rect 42476 45276 42980 45332
rect 42252 45266 42308 45276
rect 42924 45218 42980 45276
rect 43148 45330 43204 45500
rect 43148 45278 43150 45330
rect 43202 45278 43204 45330
rect 43148 45266 43204 45278
rect 43372 45332 43428 45838
rect 43820 45780 43876 45790
rect 43820 45686 43876 45724
rect 44044 45666 44100 45678
rect 44044 45614 44046 45666
rect 44098 45614 44100 45666
rect 44044 45556 44100 45614
rect 44044 45490 44100 45500
rect 43372 45266 43428 45276
rect 42924 45166 42926 45218
rect 42978 45166 42980 45218
rect 42924 45154 42980 45166
rect 43820 45106 43876 45118
rect 43820 45054 43822 45106
rect 43874 45054 43876 45106
rect 43260 44996 43316 45006
rect 43260 44902 43316 44940
rect 41356 44828 41860 44884
rect 41356 42868 41412 44828
rect 41356 42802 41412 42812
rect 43148 42868 43204 42878
rect 43204 42812 43316 42868
rect 43148 42774 43204 42812
rect 43260 42194 43316 42812
rect 43820 42756 43876 45054
rect 43820 42690 43876 42700
rect 43932 42868 43988 42878
rect 43484 42644 43540 42654
rect 43484 42550 43540 42588
rect 43820 42532 43876 42542
rect 43932 42532 43988 42812
rect 44268 42756 44324 42766
rect 44268 42662 44324 42700
rect 43260 42142 43262 42194
rect 43314 42142 43316 42194
rect 43260 42130 43316 42142
rect 43596 42530 43988 42532
rect 43596 42478 43822 42530
rect 43874 42478 43988 42530
rect 43596 42476 43988 42478
rect 43372 42084 43428 42094
rect 43596 42084 43652 42476
rect 43820 42466 43876 42476
rect 44380 42420 44436 46396
rect 44492 44996 44548 45006
rect 44492 44902 44548 44940
rect 44828 42868 44884 42878
rect 44828 42754 44884 42812
rect 44828 42702 44830 42754
rect 44882 42702 44884 42754
rect 44828 42690 44884 42702
rect 45388 42868 45444 42878
rect 45388 42754 45444 42812
rect 45388 42702 45390 42754
rect 45442 42702 45444 42754
rect 45388 42690 45444 42702
rect 45500 42642 45556 46620
rect 46060 45332 46116 45342
rect 46060 43762 46116 45276
rect 46060 43710 46062 43762
rect 46114 43710 46116 43762
rect 46060 43698 46116 43710
rect 45948 43538 46004 43550
rect 45948 43486 45950 43538
rect 46002 43486 46004 43538
rect 45948 42868 46004 43486
rect 45948 42802 46004 42812
rect 45500 42590 45502 42642
rect 45554 42590 45556 42642
rect 45500 42578 45556 42590
rect 44940 42530 44996 42542
rect 44940 42478 44942 42530
rect 44994 42478 44996 42530
rect 44940 42420 44996 42478
rect 44380 42364 44996 42420
rect 45164 42530 45220 42542
rect 45164 42478 45166 42530
rect 45218 42478 45220 42530
rect 43372 42082 43652 42084
rect 43372 42030 43374 42082
rect 43426 42030 43652 42082
rect 43372 42028 43652 42030
rect 43372 42018 43428 42028
rect 41244 41918 41246 41970
rect 41298 41918 41300 41970
rect 41244 41906 41300 41918
rect 44268 41860 44324 41870
rect 44044 41804 44268 41860
rect 41020 41692 41300 41748
rect 40348 39554 40404 39564
rect 40460 40962 40964 40964
rect 40460 40910 40574 40962
rect 40626 40910 40964 40962
rect 40460 40908 40964 40910
rect 41132 41076 41188 41086
rect 40348 37156 40404 37166
rect 40348 37062 40404 37100
rect 39788 34354 39956 34356
rect 39788 34302 39790 34354
rect 39842 34302 39956 34354
rect 39788 34300 39956 34302
rect 40012 36260 40068 36270
rect 40012 34914 40068 36204
rect 40460 36148 40516 40908
rect 40572 40898 40628 40908
rect 40796 40404 40852 40414
rect 40796 40310 40852 40348
rect 41132 40402 41188 41020
rect 41132 40350 41134 40402
rect 41186 40350 41188 40402
rect 41132 40338 41188 40350
rect 41020 40292 41076 40302
rect 40908 40290 41076 40292
rect 40908 40238 41022 40290
rect 41074 40238 41076 40290
rect 40908 40236 41076 40238
rect 40908 39844 40964 40236
rect 41020 40226 41076 40236
rect 40572 39788 40964 39844
rect 40572 39730 40628 39788
rect 40572 39678 40574 39730
rect 40626 39678 40628 39730
rect 40572 39666 40628 39678
rect 40908 39396 40964 39406
rect 40908 38052 40964 39340
rect 41244 38668 41300 41692
rect 43260 41746 43316 41758
rect 43260 41694 43262 41746
rect 43314 41694 43316 41746
rect 41804 40964 41860 40974
rect 41468 40962 41860 40964
rect 41468 40910 41806 40962
rect 41858 40910 41860 40962
rect 41468 40908 41860 40910
rect 41468 40514 41524 40908
rect 41804 40898 41860 40908
rect 42028 40628 42084 40638
rect 42028 40534 42084 40572
rect 41468 40462 41470 40514
rect 41522 40462 41524 40514
rect 41468 39844 41524 40462
rect 42364 40514 42420 40526
rect 42364 40462 42366 40514
rect 42418 40462 42420 40514
rect 42364 40292 42420 40462
rect 42364 40226 42420 40236
rect 41468 39778 41524 39788
rect 43036 39844 43092 39854
rect 41356 39620 41412 39630
rect 41804 39620 41860 39630
rect 41412 39618 41860 39620
rect 41412 39566 41806 39618
rect 41858 39566 41860 39618
rect 41412 39564 41860 39566
rect 41356 39526 41412 39564
rect 41804 39554 41860 39564
rect 43036 39060 43092 39788
rect 40908 37938 40964 37996
rect 40908 37886 40910 37938
rect 40962 37886 40964 37938
rect 40908 37874 40964 37886
rect 41020 38612 41300 38668
rect 42812 38724 42868 38762
rect 42812 38658 42868 38668
rect 40460 36082 40516 36092
rect 40908 35588 40964 35598
rect 40236 35364 40292 35374
rect 40012 34862 40014 34914
rect 40066 34862 40068 34914
rect 39788 34290 39844 34300
rect 39900 34132 39956 34142
rect 39900 34038 39956 34076
rect 39676 32622 39678 32674
rect 39730 32622 39732 32674
rect 39676 32610 39732 32622
rect 39788 33906 39844 33918
rect 39788 33854 39790 33906
rect 39842 33854 39844 33906
rect 39676 31780 39732 31790
rect 39676 31686 39732 31724
rect 39564 29708 39732 29764
rect 39452 29596 39620 29652
rect 39004 29558 39060 29596
rect 38444 29486 38446 29538
rect 38498 29486 38500 29538
rect 38220 29204 38276 29484
rect 38444 29474 38500 29486
rect 39564 29538 39620 29596
rect 39564 29486 39566 29538
rect 39618 29486 39620 29538
rect 39564 29474 39620 29486
rect 39676 29540 39732 29708
rect 39676 29474 39732 29484
rect 39004 29428 39060 29438
rect 39452 29428 39508 29438
rect 39004 29334 39060 29372
rect 39228 29426 39508 29428
rect 39228 29374 39454 29426
rect 39506 29374 39508 29426
rect 39228 29372 39508 29374
rect 38108 28868 38164 28878
rect 38220 28868 38276 29148
rect 38780 29204 38836 29214
rect 39228 29204 39284 29372
rect 39452 29362 39508 29372
rect 39564 29316 39620 29326
rect 38780 29202 39284 29204
rect 38780 29150 38782 29202
rect 38834 29150 39284 29202
rect 38780 29148 39284 29150
rect 39340 29204 39396 29214
rect 38780 29138 38836 29148
rect 39340 29110 39396 29148
rect 39564 28980 39620 29260
rect 39228 28924 39620 28980
rect 38108 28866 38276 28868
rect 38108 28814 38110 28866
rect 38162 28814 38276 28866
rect 38108 28812 38276 28814
rect 39004 28868 39060 28878
rect 38108 28802 38164 28812
rect 37772 28590 37774 28642
rect 37826 28590 37828 28642
rect 37436 28018 37492 28028
rect 37660 27860 37716 27870
rect 37660 27766 37716 27804
rect 37212 27748 37268 27758
rect 37212 27654 37268 27692
rect 37772 27076 37828 28590
rect 37772 27010 37828 27020
rect 37884 27972 37940 27982
rect 37324 26180 37380 26190
rect 37100 25618 37156 25630
rect 37100 25566 37102 25618
rect 37154 25566 37156 25618
rect 37100 25508 37156 25566
rect 37100 25442 37156 25452
rect 36988 24098 37044 24108
rect 37100 24724 37156 24734
rect 36988 22372 37044 22382
rect 37100 22372 37156 24668
rect 37324 23716 37380 26124
rect 37548 25284 37604 25294
rect 37548 25190 37604 25228
rect 37660 25060 37716 25070
rect 37660 23940 37716 25004
rect 37772 24724 37828 24734
rect 37772 24630 37828 24668
rect 37660 23846 37716 23884
rect 37324 23650 37380 23660
rect 37436 23714 37492 23726
rect 37436 23662 37438 23714
rect 37490 23662 37492 23714
rect 37436 23604 37492 23662
rect 37772 23714 37828 23726
rect 37772 23662 37774 23714
rect 37826 23662 37828 23714
rect 37772 23604 37828 23662
rect 37436 23548 37828 23604
rect 37212 23044 37268 23054
rect 37212 22950 37268 22988
rect 37100 22316 37268 22372
rect 36988 22278 37044 22316
rect 37100 22146 37156 22158
rect 37100 22094 37102 22146
rect 37154 22094 37156 22146
rect 37100 21476 37156 22094
rect 37212 21812 37268 22316
rect 37324 22260 37380 22270
rect 37324 22166 37380 22204
rect 37212 21746 37268 21756
rect 37100 21410 37156 21420
rect 36764 16706 36820 16716
rect 37100 16994 37156 17006
rect 37100 16942 37102 16994
rect 37154 16942 37156 16994
rect 37100 15874 37156 16942
rect 37100 15822 37102 15874
rect 37154 15822 37156 15874
rect 37100 15428 37156 15822
rect 37100 15362 37156 15372
rect 36988 15316 37044 15326
rect 36988 15222 37044 15260
rect 37100 12180 37156 12190
rect 37100 12086 37156 12124
rect 37436 10948 37492 23548
rect 37660 23266 37716 23278
rect 37660 23214 37662 23266
rect 37714 23214 37716 23266
rect 37548 23044 37604 23054
rect 37548 21924 37604 22988
rect 37548 20916 37604 21868
rect 37660 21476 37716 23214
rect 37884 22484 37940 27916
rect 38780 27970 38836 27982
rect 38780 27918 38782 27970
rect 38834 27918 38836 27970
rect 38780 26908 38836 27918
rect 39004 27858 39060 28812
rect 39228 28754 39284 28924
rect 39228 28702 39230 28754
rect 39282 28702 39284 28754
rect 39228 28690 39284 28702
rect 39564 28420 39620 28430
rect 39004 27806 39006 27858
rect 39058 27806 39060 27858
rect 39004 26908 39060 27806
rect 39452 28418 39620 28420
rect 39452 28366 39566 28418
rect 39618 28366 39620 28418
rect 39452 28364 39620 28366
rect 39340 27076 39396 27086
rect 39452 27076 39508 28364
rect 39564 28354 39620 28364
rect 39788 27914 39844 33854
rect 39900 32676 39956 32686
rect 40012 32676 40068 34862
rect 39956 32620 40068 32676
rect 40124 35308 40236 35364
rect 39900 32582 39956 32620
rect 39900 31780 39956 31790
rect 39900 31686 39956 31724
rect 40124 31332 40180 35308
rect 40236 35298 40292 35308
rect 40572 34916 40628 34926
rect 40796 34916 40852 34926
rect 40572 34914 40796 34916
rect 40572 34862 40574 34914
rect 40626 34862 40796 34914
rect 40572 34860 40796 34862
rect 40572 34850 40628 34860
rect 40796 34850 40852 34860
rect 40908 34690 40964 35532
rect 40908 34638 40910 34690
rect 40962 34638 40964 34690
rect 40908 34626 40964 34638
rect 41020 34130 41076 38612
rect 41244 37828 41300 37838
rect 41244 37826 41524 37828
rect 41244 37774 41246 37826
rect 41298 37774 41524 37826
rect 41244 37772 41524 37774
rect 41244 37762 41300 37772
rect 41468 34916 41524 37772
rect 42364 37380 42420 37390
rect 42028 37044 42084 37054
rect 41580 35588 41636 35598
rect 41580 35586 41748 35588
rect 41580 35534 41582 35586
rect 41634 35534 41748 35586
rect 41580 35532 41748 35534
rect 41580 35522 41636 35532
rect 41580 34916 41636 34926
rect 41020 34078 41022 34130
rect 41074 34078 41076 34130
rect 41020 33460 41076 34078
rect 40684 33122 40740 33134
rect 40684 33070 40686 33122
rect 40738 33070 40740 33122
rect 40460 32676 40516 32686
rect 40460 32582 40516 32620
rect 40684 32564 40740 33070
rect 40908 32564 40964 32574
rect 40684 32562 40964 32564
rect 40684 32510 40910 32562
rect 40962 32510 40964 32562
rect 40684 32508 40964 32510
rect 40236 32004 40292 32014
rect 40236 31666 40292 31948
rect 40908 32004 40964 32508
rect 40908 31938 40964 31948
rect 40236 31614 40238 31666
rect 40290 31614 40292 31666
rect 40236 31602 40292 31614
rect 40348 31780 40404 31790
rect 40348 31444 40404 31724
rect 40012 31276 40180 31332
rect 40236 31388 40404 31444
rect 40684 31778 40740 31790
rect 40684 31726 40686 31778
rect 40738 31726 40740 31778
rect 39900 29426 39956 29438
rect 39900 29374 39902 29426
rect 39954 29374 39956 29426
rect 39900 28642 39956 29374
rect 39900 28590 39902 28642
rect 39954 28590 39956 28642
rect 39900 28578 39956 28590
rect 40012 28084 40068 31276
rect 40236 29538 40292 31388
rect 40236 29486 40238 29538
rect 40290 29486 40292 29538
rect 40124 29428 40180 29438
rect 40236 29428 40292 29486
rect 40348 29540 40404 29550
rect 40348 29446 40404 29484
rect 40124 29426 40292 29428
rect 40124 29374 40126 29426
rect 40178 29374 40292 29426
rect 40124 29372 40292 29374
rect 40124 29362 40180 29372
rect 40236 29316 40292 29372
rect 40684 29428 40740 31726
rect 41020 31780 41076 33404
rect 41020 31714 41076 31724
rect 41132 34860 41468 34916
rect 41524 34914 41636 34916
rect 41524 34862 41582 34914
rect 41634 34862 41636 34914
rect 41524 34860 41636 34862
rect 41132 32788 41188 34860
rect 41468 34822 41524 34860
rect 41580 34850 41636 34860
rect 41244 34692 41300 34702
rect 41692 34692 41748 35532
rect 41244 34690 41748 34692
rect 41244 34638 41246 34690
rect 41298 34638 41748 34690
rect 41244 34636 41748 34638
rect 41916 34692 41972 34702
rect 41244 34626 41300 34636
rect 41356 34018 41412 34636
rect 41916 34598 41972 34636
rect 41356 33966 41358 34018
rect 41410 33966 41412 34018
rect 41244 32788 41300 32798
rect 41132 32786 41300 32788
rect 41132 32734 41246 32786
rect 41298 32734 41300 32786
rect 41132 32732 41300 32734
rect 41132 31778 41188 32732
rect 41244 32722 41300 32732
rect 41132 31726 41134 31778
rect 41186 31726 41188 31778
rect 41132 31714 41188 31726
rect 41356 31556 41412 33966
rect 42028 33908 42084 36988
rect 42364 35588 42420 37324
rect 42700 37156 42756 37166
rect 43036 37156 43092 39004
rect 43260 37378 43316 41694
rect 44044 40626 44100 41804
rect 44268 41794 44324 41804
rect 44940 41860 44996 41870
rect 44996 41804 45108 41860
rect 44940 41794 44996 41804
rect 44044 40574 44046 40626
rect 44098 40574 44100 40626
rect 44044 40562 44100 40574
rect 44268 41076 44324 41086
rect 44268 40626 44324 41020
rect 44268 40574 44270 40626
rect 44322 40574 44324 40626
rect 44268 40562 44324 40574
rect 43708 40516 43764 40526
rect 43708 40422 43764 40460
rect 44492 40516 44548 40526
rect 43932 40402 43988 40414
rect 43932 40350 43934 40402
rect 43986 40350 43988 40402
rect 43932 40292 43988 40350
rect 44492 40404 44548 40460
rect 44492 40402 44884 40404
rect 44492 40350 44494 40402
rect 44546 40350 44884 40402
rect 44492 40348 44884 40350
rect 44492 40338 44548 40348
rect 43988 40236 44100 40292
rect 43932 40226 43988 40236
rect 44044 39620 44100 40236
rect 44044 39618 44324 39620
rect 44044 39566 44046 39618
rect 44098 39566 44324 39618
rect 44044 39564 44324 39566
rect 44044 39554 44100 39564
rect 44268 39508 44324 39564
rect 44156 39394 44212 39406
rect 44156 39342 44158 39394
rect 44210 39342 44212 39394
rect 44156 38948 44212 39342
rect 43932 38892 44212 38948
rect 43932 38724 43988 38892
rect 44268 38836 44324 39452
rect 44716 39618 44772 39630
rect 44716 39566 44718 39618
rect 44770 39566 44772 39618
rect 44380 39396 44436 39406
rect 44716 39396 44772 39566
rect 44380 39394 44772 39396
rect 44380 39342 44382 39394
rect 44434 39342 44772 39394
rect 44380 39340 44772 39342
rect 44380 39330 44436 39340
rect 43820 37380 43876 37390
rect 43260 37326 43262 37378
rect 43314 37326 43316 37378
rect 43260 37314 43316 37326
rect 43708 37378 43876 37380
rect 43708 37326 43822 37378
rect 43874 37326 43876 37378
rect 43708 37324 43876 37326
rect 43148 37266 43204 37278
rect 43148 37214 43150 37266
rect 43202 37214 43204 37266
rect 43148 37156 43204 37214
rect 43708 37266 43764 37324
rect 43820 37314 43876 37324
rect 43708 37214 43710 37266
rect 43762 37214 43764 37266
rect 43708 37202 43764 37214
rect 42700 37154 43204 37156
rect 42700 37102 42702 37154
rect 42754 37102 43204 37154
rect 42700 37100 43204 37102
rect 42700 37090 42756 37100
rect 42364 35586 42644 35588
rect 42364 35534 42366 35586
rect 42418 35534 42644 35586
rect 42364 35532 42644 35534
rect 42364 35522 42420 35532
rect 42588 34802 42644 35532
rect 42812 35028 42868 35038
rect 42588 34750 42590 34802
rect 42642 34750 42644 34802
rect 42588 34738 42644 34750
rect 42700 34802 42756 34814
rect 42700 34750 42702 34802
rect 42754 34750 42756 34802
rect 42364 34690 42420 34702
rect 42364 34638 42366 34690
rect 42418 34638 42420 34690
rect 42140 34242 42196 34254
rect 42140 34190 42142 34242
rect 42194 34190 42196 34242
rect 42140 34132 42196 34190
rect 42140 34066 42196 34076
rect 42028 33852 42196 33908
rect 41468 33460 41524 33470
rect 41692 33460 41748 33470
rect 41524 33458 41748 33460
rect 41524 33406 41694 33458
rect 41746 33406 41748 33458
rect 41524 33404 41748 33406
rect 41468 33394 41524 33404
rect 41692 33394 41748 33404
rect 41804 33460 41860 33470
rect 40236 29260 40628 29316
rect 40572 28866 40628 29260
rect 40572 28814 40574 28866
rect 40626 28814 40628 28866
rect 40572 28754 40628 28814
rect 40572 28702 40574 28754
rect 40626 28702 40628 28754
rect 40572 28690 40628 28702
rect 40236 28308 40292 28318
rect 40012 28028 40180 28084
rect 39788 27862 39790 27914
rect 39842 27862 39844 27914
rect 39788 27850 39844 27862
rect 40012 27860 40068 27870
rect 39900 27858 40068 27860
rect 39900 27806 40014 27858
rect 40066 27806 40068 27858
rect 39900 27804 40068 27806
rect 39788 27636 39844 27646
rect 39788 27188 39844 27580
rect 39788 27094 39844 27132
rect 39340 27074 39508 27076
rect 39340 27022 39342 27074
rect 39394 27022 39508 27074
rect 39340 27020 39508 27022
rect 39340 27010 39396 27020
rect 37996 26852 38052 26862
rect 37996 25844 38052 26796
rect 37996 25618 38052 25788
rect 38668 26852 38836 26908
rect 38892 26852 39060 26908
rect 38668 25732 38724 26852
rect 38892 26404 38948 26852
rect 39452 26740 39508 27020
rect 39900 26964 39956 27804
rect 40012 27794 40068 27804
rect 40124 26908 40180 28028
rect 40236 27970 40292 28252
rect 40236 27918 40238 27970
rect 40290 27918 40292 27970
rect 40236 27906 40292 27918
rect 39900 26898 39956 26908
rect 39452 26674 39508 26684
rect 40012 26852 40180 26908
rect 40236 26962 40292 26974
rect 40236 26910 40238 26962
rect 40290 26910 40292 26962
rect 38892 26402 39060 26404
rect 38892 26350 38894 26402
rect 38946 26350 39060 26402
rect 38892 26348 39060 26350
rect 38892 26338 38948 26348
rect 38780 26292 38836 26302
rect 38780 26198 38836 26236
rect 38892 26068 38948 26078
rect 38892 25974 38948 26012
rect 39004 25844 39060 26348
rect 39676 26068 39732 26078
rect 38668 25666 38724 25676
rect 38892 25788 39060 25844
rect 39340 25844 39396 25854
rect 37996 25566 37998 25618
rect 38050 25566 38052 25618
rect 37996 25554 38052 25566
rect 38108 25508 38164 25518
rect 37996 23828 38052 23838
rect 37996 23734 38052 23772
rect 38108 23154 38164 25452
rect 38556 25284 38612 25294
rect 38556 25190 38612 25228
rect 38556 24724 38612 24734
rect 38556 24630 38612 24668
rect 38780 23828 38836 23838
rect 38780 23734 38836 23772
rect 38892 23826 38948 25788
rect 38892 23774 38894 23826
rect 38946 23774 38948 23826
rect 38892 23762 38948 23774
rect 39004 25506 39060 25518
rect 39004 25454 39006 25506
rect 39058 25454 39060 25506
rect 38108 23102 38110 23154
rect 38162 23102 38164 23154
rect 38108 23090 38164 23102
rect 38444 23154 38500 23166
rect 38444 23102 38446 23154
rect 38498 23102 38500 23154
rect 38444 23044 38500 23102
rect 38444 22978 38500 22988
rect 37996 22484 38052 22494
rect 38668 22484 38724 22494
rect 37884 22482 38052 22484
rect 37884 22430 37998 22482
rect 38050 22430 38052 22482
rect 37884 22428 38052 22430
rect 37996 21700 38052 22428
rect 38556 22482 38724 22484
rect 38556 22430 38670 22482
rect 38722 22430 38724 22482
rect 38556 22428 38724 22430
rect 38556 21812 38612 22428
rect 38668 22418 38724 22428
rect 38556 21718 38612 21756
rect 37996 21634 38052 21644
rect 37660 21410 37716 21420
rect 38108 21476 38164 21486
rect 37548 20850 37604 20860
rect 38108 20188 38164 21420
rect 37660 20132 38164 20188
rect 37660 17666 37716 20132
rect 39004 19684 39060 25454
rect 39340 25396 39396 25788
rect 39340 25302 39396 25340
rect 39676 25394 39732 26012
rect 39676 25342 39678 25394
rect 39730 25342 39732 25394
rect 39676 25330 39732 25342
rect 39788 25506 39844 25518
rect 39788 25454 39790 25506
rect 39842 25454 39844 25506
rect 39452 24948 39508 24958
rect 39228 24834 39284 24846
rect 39228 24782 39230 24834
rect 39282 24782 39284 24834
rect 39116 23940 39172 23950
rect 39228 23940 39284 24782
rect 39452 24724 39508 24892
rect 39788 24948 39844 25454
rect 39788 24882 39844 24892
rect 39900 25396 39956 25406
rect 39900 24834 39956 25340
rect 40012 25282 40068 26852
rect 40012 25230 40014 25282
rect 40066 25230 40068 25282
rect 40012 25218 40068 25230
rect 40124 26740 40180 26750
rect 40236 26740 40292 26910
rect 40180 26684 40292 26740
rect 39900 24782 39902 24834
rect 39954 24782 39956 24834
rect 39900 24770 39956 24782
rect 39116 23938 39284 23940
rect 39116 23886 39118 23938
rect 39170 23886 39284 23938
rect 39116 23884 39284 23886
rect 39340 24722 39508 24724
rect 39340 24670 39454 24722
rect 39506 24670 39508 24722
rect 39340 24668 39508 24670
rect 39116 23874 39172 23884
rect 39340 23492 39396 24668
rect 39452 24658 39508 24668
rect 40012 24722 40068 24734
rect 40012 24670 40014 24722
rect 40066 24670 40068 24722
rect 39676 24612 39732 24622
rect 39564 23940 39620 23950
rect 39228 23436 39396 23492
rect 39452 23492 39508 23502
rect 39228 23154 39284 23436
rect 39340 23268 39396 23278
rect 39452 23268 39508 23436
rect 39340 23266 39508 23268
rect 39340 23214 39342 23266
rect 39394 23214 39508 23266
rect 39340 23212 39508 23214
rect 39564 23266 39620 23884
rect 39564 23214 39566 23266
rect 39618 23214 39620 23266
rect 39340 23202 39396 23212
rect 39564 23202 39620 23214
rect 39228 23102 39230 23154
rect 39282 23102 39284 23154
rect 39228 22372 39284 23102
rect 39228 22306 39284 22316
rect 39228 21700 39284 21710
rect 39228 20914 39284 21644
rect 39228 20862 39230 20914
rect 39282 20862 39284 20914
rect 39228 20850 39284 20862
rect 39564 21474 39620 21486
rect 39564 21422 39566 21474
rect 39618 21422 39620 21474
rect 39564 20580 39620 21422
rect 39564 20514 39620 20524
rect 39004 19618 39060 19628
rect 39676 19572 39732 24556
rect 40012 24500 40068 24670
rect 40012 23548 40068 24444
rect 39900 23492 40068 23548
rect 39788 19796 39844 19806
rect 39788 19702 39844 19740
rect 39788 19572 39844 19582
rect 39676 19516 39788 19572
rect 39788 19506 39844 19516
rect 38444 19460 38500 19470
rect 38444 19366 38500 19404
rect 39452 19346 39508 19358
rect 39452 19294 39454 19346
rect 39506 19294 39508 19346
rect 38668 19124 38724 19134
rect 39116 19124 39172 19134
rect 38668 19122 39172 19124
rect 38668 19070 38670 19122
rect 38722 19070 39118 19122
rect 39170 19070 39172 19122
rect 38668 19068 39172 19070
rect 38668 19058 38724 19068
rect 39116 19058 39172 19068
rect 38556 19010 38612 19022
rect 38556 18958 38558 19010
rect 38610 18958 38612 19010
rect 38332 18674 38388 18686
rect 38332 18622 38334 18674
rect 38386 18622 38388 18674
rect 38332 18564 38388 18622
rect 38332 18498 38388 18508
rect 38556 17780 38612 18958
rect 38892 18452 38948 18462
rect 38892 18358 38948 18396
rect 38556 17714 38612 17724
rect 37660 17614 37662 17666
rect 37714 17614 37716 17666
rect 37660 17602 37716 17614
rect 37996 17666 38052 17678
rect 37996 17614 37998 17666
rect 38050 17614 38052 17666
rect 37884 17444 37940 17454
rect 37548 16884 37604 16894
rect 37548 16882 37716 16884
rect 37548 16830 37550 16882
rect 37602 16830 37716 16882
rect 37548 16828 37716 16830
rect 37548 16818 37604 16828
rect 37436 10882 37492 10892
rect 37660 15428 37716 16828
rect 37884 16882 37940 17388
rect 37884 16830 37886 16882
rect 37938 16830 37940 16882
rect 37884 16818 37940 16830
rect 37996 16098 38052 17614
rect 38108 17668 38164 17678
rect 38108 17574 38164 17612
rect 39116 17666 39172 17678
rect 39116 17614 39118 17666
rect 39170 17614 39172 17666
rect 38556 17556 38612 17566
rect 38612 17500 39060 17556
rect 38556 17462 38612 17500
rect 37996 16046 37998 16098
rect 38050 16046 38052 16098
rect 37772 15876 37828 15886
rect 37772 15782 37828 15820
rect 37996 15876 38052 16046
rect 38108 17106 38164 17118
rect 38108 17054 38110 17106
rect 38162 17054 38164 17106
rect 38108 15988 38164 17054
rect 38332 17106 38388 17118
rect 38332 17054 38334 17106
rect 38386 17054 38388 17106
rect 38220 16436 38276 16446
rect 38220 15988 38276 16380
rect 38332 16212 38388 17054
rect 39004 17106 39060 17500
rect 39004 17054 39006 17106
rect 39058 17054 39060 17106
rect 39004 17042 39060 17054
rect 38668 16324 38724 16334
rect 38556 16212 38612 16222
rect 38332 16156 38556 16212
rect 38556 16098 38612 16156
rect 38556 16046 38558 16098
rect 38610 16046 38612 16098
rect 38556 16034 38612 16046
rect 38668 16098 38724 16268
rect 38668 16046 38670 16098
rect 38722 16046 38724 16098
rect 38332 15988 38388 15998
rect 38220 15986 38388 15988
rect 38220 15934 38334 15986
rect 38386 15934 38388 15986
rect 38220 15932 38388 15934
rect 38108 15922 38164 15932
rect 37996 15810 38052 15820
rect 37660 15372 38052 15428
rect 37660 10052 37716 15372
rect 37996 15314 38052 15372
rect 37996 15262 37998 15314
rect 38050 15262 38052 15314
rect 37996 15250 38052 15262
rect 38332 15204 38388 15932
rect 38668 15652 38724 16046
rect 39116 15764 39172 17614
rect 39452 16436 39508 19294
rect 39788 19236 39844 19246
rect 39900 19236 39956 23492
rect 40012 23156 40068 23166
rect 40012 23062 40068 23100
rect 40012 22372 40068 22382
rect 40012 21698 40068 22316
rect 40012 21646 40014 21698
rect 40066 21646 40068 21698
rect 40012 21634 40068 21646
rect 40124 20244 40180 26684
rect 40236 25172 40292 25182
rect 40236 24610 40292 25116
rect 40236 24558 40238 24610
rect 40290 24558 40292 24610
rect 40236 24546 40292 24558
rect 40348 22370 40404 22382
rect 40348 22318 40350 22370
rect 40402 22318 40404 22370
rect 40348 21700 40404 22318
rect 40348 21634 40404 21644
rect 40460 22148 40516 22158
rect 40124 20178 40180 20188
rect 40236 21588 40292 21598
rect 40124 20020 40180 20030
rect 40236 20020 40292 21532
rect 40124 20018 40292 20020
rect 40124 19966 40126 20018
rect 40178 19966 40292 20018
rect 40124 19964 40292 19966
rect 40348 20020 40404 20030
rect 40460 20020 40516 22092
rect 40348 20018 40516 20020
rect 40348 19966 40350 20018
rect 40402 19966 40516 20018
rect 40348 19964 40516 19966
rect 40124 19954 40180 19964
rect 40348 19954 40404 19964
rect 39788 19234 39956 19236
rect 39788 19182 39790 19234
rect 39842 19182 39956 19234
rect 39788 19180 39956 19182
rect 39788 19170 39844 19180
rect 40348 18452 40404 18462
rect 39452 16370 39508 16380
rect 39564 17780 39620 17790
rect 39564 15988 39620 17724
rect 40012 17442 40068 17454
rect 40012 17390 40014 17442
rect 40066 17390 40068 17442
rect 40012 16098 40068 17390
rect 40012 16046 40014 16098
rect 40066 16046 40068 16098
rect 40012 16034 40068 16046
rect 39676 15988 39732 15998
rect 39564 15986 39732 15988
rect 39564 15934 39678 15986
rect 39730 15934 39732 15986
rect 39564 15932 39732 15934
rect 39676 15922 39732 15932
rect 38668 15586 38724 15596
rect 38780 15708 39172 15764
rect 38332 15138 38388 15148
rect 38444 15428 38500 15438
rect 38444 15202 38500 15372
rect 38444 15150 38446 15202
rect 38498 15150 38500 15202
rect 38444 15138 38500 15150
rect 38780 14980 38836 15708
rect 39564 15540 39620 15550
rect 38668 14532 38724 14542
rect 38780 14532 38836 14924
rect 38892 15090 38948 15102
rect 38892 15038 38894 15090
rect 38946 15038 38948 15090
rect 38892 14868 38948 15038
rect 38892 14812 39284 14868
rect 38668 14530 38836 14532
rect 38668 14478 38670 14530
rect 38722 14478 38836 14530
rect 38668 14476 38836 14478
rect 38892 14644 38948 14654
rect 38892 14530 38948 14588
rect 38892 14478 38894 14530
rect 38946 14478 38948 14530
rect 38668 14466 38724 14476
rect 38892 14466 38948 14478
rect 38108 14420 38164 14430
rect 39116 14420 39172 14430
rect 38108 13188 38164 14364
rect 38108 12962 38164 13132
rect 39004 14418 39172 14420
rect 39004 14366 39118 14418
rect 39170 14366 39172 14418
rect 39004 14364 39172 14366
rect 38108 12910 38110 12962
rect 38162 12910 38164 12962
rect 38108 12898 38164 12910
rect 38332 12964 38388 12974
rect 38332 12870 38388 12908
rect 38780 12964 38836 12974
rect 39004 12964 39060 14364
rect 39116 14354 39172 14364
rect 39228 13300 39284 14812
rect 39228 13234 39284 13244
rect 38780 12962 39060 12964
rect 38780 12910 38782 12962
rect 38834 12910 39060 12962
rect 38780 12908 39060 12910
rect 38780 12898 38836 12908
rect 37772 12740 37828 12750
rect 37772 10500 37828 12684
rect 38444 12738 38500 12750
rect 38444 12686 38446 12738
rect 38498 12686 38500 12738
rect 37884 12068 37940 12078
rect 37884 12066 38164 12068
rect 37884 12014 37886 12066
rect 37938 12014 38164 12066
rect 37884 12012 38164 12014
rect 37884 12002 37940 12012
rect 38108 11618 38164 12012
rect 38108 11566 38110 11618
rect 38162 11566 38164 11618
rect 38108 11554 38164 11566
rect 38220 11844 38276 11854
rect 38220 11282 38276 11788
rect 38444 11618 38500 12686
rect 38556 12740 38612 12750
rect 38556 12646 38612 12684
rect 38444 11566 38446 11618
rect 38498 11566 38500 11618
rect 38444 11554 38500 11566
rect 38220 11230 38222 11282
rect 38274 11230 38276 11282
rect 38220 11218 38276 11230
rect 39452 10836 39508 10846
rect 39564 10836 39620 15484
rect 39788 15428 39844 15438
rect 39340 10834 39620 10836
rect 39340 10782 39454 10834
rect 39506 10782 39620 10834
rect 39340 10780 39620 10782
rect 39676 14308 39732 14318
rect 39676 13970 39732 14252
rect 39676 13918 39678 13970
rect 39730 13918 39732 13970
rect 37772 10444 38052 10500
rect 37660 9986 37716 9996
rect 37100 9826 37156 9838
rect 37100 9774 37102 9826
rect 37154 9774 37156 9826
rect 37100 9604 37156 9774
rect 37996 9714 38052 10444
rect 39228 10388 39284 10398
rect 39004 10386 39284 10388
rect 39004 10334 39230 10386
rect 39282 10334 39284 10386
rect 39004 10332 39284 10334
rect 38220 9828 38276 9838
rect 38220 9734 38276 9772
rect 38668 9828 38724 9838
rect 38668 9734 38724 9772
rect 39004 9826 39060 10332
rect 39228 10322 39284 10332
rect 39004 9774 39006 9826
rect 39058 9774 39060 9826
rect 39004 9762 39060 9774
rect 39228 9828 39284 9838
rect 39340 9828 39396 10780
rect 39452 10770 39508 10780
rect 39228 9826 39396 9828
rect 39228 9774 39230 9826
rect 39282 9774 39396 9826
rect 39228 9772 39396 9774
rect 39676 9828 39732 13918
rect 39788 12964 39844 15372
rect 39900 15090 39956 15102
rect 39900 15038 39902 15090
rect 39954 15038 39956 15090
rect 39900 14980 39956 15038
rect 39900 14914 39956 14924
rect 40236 14980 40292 14990
rect 40012 14196 40068 14206
rect 40012 13970 40068 14140
rect 40012 13918 40014 13970
rect 40066 13918 40068 13970
rect 40012 13906 40068 13918
rect 40012 12964 40068 12974
rect 39788 12908 40012 12964
rect 37996 9662 37998 9714
rect 38050 9662 38052 9714
rect 37100 9538 37156 9548
rect 37324 9602 37380 9614
rect 37324 9550 37326 9602
rect 37378 9550 37380 9602
rect 35980 8372 36148 8428
rect 36428 8372 36708 8428
rect 35980 7698 36036 8372
rect 35980 7646 35982 7698
rect 36034 7646 36036 7698
rect 35980 7634 36036 7646
rect 35812 7420 36148 7476
rect 35756 7410 35812 7420
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 33292 6916 33348 6926
rect 32284 6638 32286 6690
rect 32338 6638 32340 6690
rect 32284 6626 32340 6638
rect 32956 6690 33012 6702
rect 32956 6638 32958 6690
rect 33010 6638 33012 6690
rect 31724 6578 31780 6590
rect 31948 6580 32004 6590
rect 31724 6526 31726 6578
rect 31778 6526 31780 6578
rect 31724 6132 31780 6526
rect 31724 6066 31780 6076
rect 31836 6578 32004 6580
rect 31836 6526 31950 6578
rect 32002 6526 32004 6578
rect 31836 6524 32004 6526
rect 31500 5348 31556 5358
rect 31836 5348 31892 6524
rect 31948 6514 32004 6524
rect 32508 6580 32564 6590
rect 32508 6466 32564 6524
rect 32508 6414 32510 6466
rect 32562 6414 32564 6466
rect 32508 6402 32564 6414
rect 31556 5292 31892 5348
rect 31500 5254 31556 5292
rect 30604 5236 30660 5246
rect 30436 5234 30660 5236
rect 30436 5182 30606 5234
rect 30658 5182 30660 5234
rect 30436 5180 30660 5182
rect 30380 5142 30436 5180
rect 30604 5170 30660 5180
rect 32956 5236 33012 6638
rect 33068 6132 33124 6142
rect 33068 6038 33124 6076
rect 33292 6130 33348 6860
rect 35756 6802 35812 6814
rect 35756 6750 35758 6802
rect 35810 6750 35812 6802
rect 33628 6580 33684 6590
rect 35756 6580 35812 6750
rect 36092 6802 36148 7420
rect 36092 6750 36094 6802
rect 36146 6750 36148 6802
rect 36092 6738 36148 6750
rect 36204 6804 36260 6814
rect 36204 6710 36260 6748
rect 36428 6690 36484 8372
rect 37324 8260 37380 9550
rect 37660 9604 37716 9614
rect 37660 9266 37716 9548
rect 37996 9268 38052 9662
rect 37660 9214 37662 9266
rect 37714 9214 37716 9266
rect 37660 9202 37716 9214
rect 37772 9212 37996 9268
rect 36428 6638 36430 6690
rect 36482 6638 36484 6690
rect 36428 6580 36484 6638
rect 35756 6524 36484 6580
rect 36876 8204 37324 8260
rect 33628 6486 33684 6524
rect 33292 6078 33294 6130
rect 33346 6078 33348 6130
rect 33292 6066 33348 6078
rect 35868 6130 35924 6524
rect 36876 6132 36932 8204
rect 37324 8194 37380 8204
rect 37548 7588 37604 7598
rect 37436 7362 37492 7374
rect 37436 7310 37438 7362
rect 37490 7310 37492 7362
rect 37436 6580 37492 7310
rect 37548 6916 37604 7532
rect 37548 6914 37716 6916
rect 37548 6862 37550 6914
rect 37602 6862 37716 6914
rect 37548 6860 37716 6862
rect 37548 6850 37604 6860
rect 37436 6132 37492 6524
rect 35868 6078 35870 6130
rect 35922 6078 35924 6130
rect 35868 6066 35924 6078
rect 36316 6130 36932 6132
rect 36316 6078 36878 6130
rect 36930 6078 36932 6130
rect 36316 6076 36932 6078
rect 36204 6018 36260 6030
rect 36204 5966 36206 6018
rect 36258 5966 36260 6018
rect 33740 5908 33796 5918
rect 33740 5814 33796 5852
rect 35980 5908 36036 5918
rect 36204 5908 36260 5966
rect 36316 6018 36372 6076
rect 36876 6066 36932 6076
rect 37100 6076 37492 6132
rect 37660 6132 37716 6860
rect 37772 6914 37828 9212
rect 37996 9202 38052 9212
rect 38892 9602 38948 9614
rect 38892 9550 38894 9602
rect 38946 9550 38948 9602
rect 38332 8146 38388 8158
rect 38332 8094 38334 8146
rect 38386 8094 38388 8146
rect 37996 8036 38052 8046
rect 37996 7942 38052 7980
rect 38220 8034 38276 8046
rect 38220 7982 38222 8034
rect 38274 7982 38276 8034
rect 37772 6862 37774 6914
rect 37826 6862 37828 6914
rect 37772 6850 37828 6862
rect 38220 6914 38276 7982
rect 38332 7812 38388 8094
rect 38332 7746 38388 7756
rect 38220 6862 38222 6914
rect 38274 6862 38276 6914
rect 38220 6850 38276 6862
rect 38780 7364 38836 7374
rect 38332 6802 38388 6814
rect 38332 6750 38334 6802
rect 38386 6750 38388 6802
rect 38220 6692 38276 6702
rect 38220 6598 38276 6636
rect 38332 6580 38388 6750
rect 38780 6802 38836 7308
rect 38780 6750 38782 6802
rect 38834 6750 38836 6802
rect 38780 6692 38836 6750
rect 38780 6626 38836 6636
rect 38332 6514 38388 6524
rect 38892 6244 38948 9550
rect 39228 9604 39284 9772
rect 39228 9538 39284 9548
rect 39676 8818 39732 9772
rect 39676 8766 39678 8818
rect 39730 8766 39732 8818
rect 39676 8754 39732 8766
rect 39788 12740 39844 12750
rect 39564 8036 39620 8046
rect 39564 7586 39620 7980
rect 39564 7534 39566 7586
rect 39618 7534 39620 7586
rect 39564 7522 39620 7534
rect 39228 6580 39284 6590
rect 39228 6486 39284 6524
rect 38780 6188 38948 6244
rect 37660 6076 38388 6132
rect 36316 5966 36318 6018
rect 36370 5966 36372 6018
rect 36316 5954 36372 5966
rect 35980 5814 36036 5852
rect 36092 5852 36204 5908
rect 30156 5070 30158 5122
rect 30210 5070 30212 5122
rect 30156 5058 30212 5070
rect 31612 5122 31668 5134
rect 31612 5070 31614 5122
rect 31666 5070 31668 5122
rect 28140 4958 28142 5010
rect 28194 4958 28196 5010
rect 28140 4946 28196 4958
rect 28364 5012 28420 5022
rect 28364 4918 28420 4956
rect 29148 5010 29204 5022
rect 29148 4958 29150 5010
rect 29202 4958 29204 5010
rect 28140 4228 28196 4238
rect 28028 4226 28196 4228
rect 28028 4174 28142 4226
rect 28194 4174 28196 4226
rect 28028 4172 28196 4174
rect 28140 4162 28196 4172
rect 28812 4228 28868 4238
rect 29148 4228 29204 4958
rect 31612 5012 31668 5070
rect 31612 4946 31668 4956
rect 32172 5012 32228 5022
rect 29708 4898 29764 4910
rect 29708 4846 29710 4898
rect 29762 4846 29764 4898
rect 29708 4564 29764 4846
rect 29708 4508 30100 4564
rect 30044 4450 30100 4508
rect 30044 4398 30046 4450
rect 30098 4398 30100 4450
rect 30044 4386 30100 4398
rect 28868 4172 29204 4228
rect 29260 4340 29316 4350
rect 28812 4134 28868 4172
rect 25004 3614 25006 3666
rect 25058 3614 25060 3666
rect 25004 3602 25060 3614
rect 29036 3668 29092 3678
rect 29260 3668 29316 4284
rect 32172 4226 32228 4956
rect 32956 4340 33012 5180
rect 33180 5794 33236 5806
rect 33180 5742 33182 5794
rect 33234 5742 33236 5794
rect 33180 4452 33236 5742
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 36092 4562 36148 5852
rect 36204 5842 36260 5852
rect 36428 5236 36484 5246
rect 36428 5142 36484 5180
rect 36876 5236 36932 5246
rect 36876 5124 36932 5180
rect 36876 5068 37044 5124
rect 36092 4510 36094 4562
rect 36146 4510 36148 4562
rect 36092 4498 36148 4510
rect 36988 4564 37044 5068
rect 37100 4676 37156 6076
rect 37212 5908 37268 5918
rect 37212 5814 37268 5852
rect 38332 5346 38388 6076
rect 38332 5294 38334 5346
rect 38386 5294 38388 5346
rect 38332 5282 38388 5294
rect 37212 5124 37268 5134
rect 37996 5124 38052 5134
rect 37212 5122 38052 5124
rect 37212 5070 37214 5122
rect 37266 5070 37998 5122
rect 38050 5070 38052 5122
rect 37212 5068 38052 5070
rect 37212 5058 37268 5068
rect 37996 5058 38052 5068
rect 38780 5122 38836 6188
rect 38780 5070 38782 5122
rect 38834 5070 38836 5122
rect 38780 5058 38836 5070
rect 39788 5124 39844 12684
rect 40012 12066 40068 12908
rect 40012 12014 40014 12066
rect 40066 12014 40068 12066
rect 40012 12002 40068 12014
rect 40236 11732 40292 14924
rect 40348 12404 40404 18396
rect 40684 18228 40740 29372
rect 40796 31500 41412 31556
rect 41804 33012 41860 33404
rect 40796 25620 40852 31500
rect 40908 30324 40964 30334
rect 40908 26180 40964 30268
rect 41356 30210 41412 30222
rect 41356 30158 41358 30210
rect 41410 30158 41412 30210
rect 41132 29988 41188 29998
rect 41132 29894 41188 29932
rect 41244 29540 41300 29550
rect 41356 29540 41412 30158
rect 41804 29540 41860 32956
rect 42028 29988 42084 29998
rect 42028 29894 42084 29932
rect 42028 29764 42084 29774
rect 42140 29764 42196 33852
rect 42364 31780 42420 34638
rect 42476 34130 42532 34142
rect 42476 34078 42478 34130
rect 42530 34078 42532 34130
rect 42476 33572 42532 34078
rect 42700 34132 42756 34750
rect 42700 34066 42756 34076
rect 42812 34130 42868 34972
rect 43148 34692 43204 37100
rect 43484 37154 43540 37166
rect 43484 37102 43486 37154
rect 43538 37102 43540 37154
rect 43484 35812 43540 37102
rect 43932 36708 43988 38668
rect 44044 38780 44324 38836
rect 44044 38668 44100 38780
rect 44044 38612 44212 38668
rect 44044 37380 44100 37390
rect 44044 37286 44100 37324
rect 44156 37378 44212 38612
rect 44268 38164 44324 38174
rect 44828 38164 44884 40348
rect 44940 39394 44996 39406
rect 44940 39342 44942 39394
rect 44994 39342 44996 39394
rect 44940 38946 44996 39342
rect 44940 38894 44942 38946
rect 44994 38894 44996 38946
rect 44940 38882 44996 38894
rect 44268 38162 44884 38164
rect 44268 38110 44270 38162
rect 44322 38110 44884 38162
rect 44268 38108 44884 38110
rect 44268 38098 44324 38108
rect 44828 38050 44884 38108
rect 44828 37998 44830 38050
rect 44882 37998 44884 38050
rect 44828 37986 44884 37998
rect 44156 37326 44158 37378
rect 44210 37326 44212 37378
rect 44156 37314 44212 37326
rect 43484 35746 43540 35756
rect 43820 36652 43988 36708
rect 43820 34802 43876 36652
rect 44044 36372 44100 36382
rect 43932 35028 43988 35038
rect 43932 34914 43988 34972
rect 43932 34862 43934 34914
rect 43986 34862 43988 34914
rect 43932 34850 43988 34862
rect 43820 34750 43822 34802
rect 43874 34750 43876 34802
rect 43820 34738 43876 34750
rect 43596 34692 43652 34702
rect 43148 34626 43204 34636
rect 43484 34690 43652 34692
rect 43484 34638 43598 34690
rect 43650 34638 43652 34690
rect 43484 34636 43652 34638
rect 42812 34078 42814 34130
rect 42866 34078 42868 34130
rect 42812 34066 42868 34078
rect 43372 34130 43428 34142
rect 43372 34078 43374 34130
rect 43426 34078 43428 34130
rect 42476 33506 42532 33516
rect 43372 33572 43428 34078
rect 43372 33012 43428 33516
rect 43372 32946 43428 32956
rect 43372 32788 43428 32798
rect 43484 32788 43540 34636
rect 43596 34626 43652 34636
rect 44044 34580 44100 36316
rect 44492 35812 44548 35822
rect 44492 35718 44548 35756
rect 44828 35028 44884 35038
rect 44828 34914 44884 34972
rect 44828 34862 44830 34914
rect 44882 34862 44884 34914
rect 44828 34850 44884 34862
rect 44940 34804 44996 34814
rect 45052 34804 45108 41804
rect 45164 39618 45220 42478
rect 45724 42530 45780 42542
rect 45724 42478 45726 42530
rect 45778 42478 45780 42530
rect 45276 41860 45332 41870
rect 45276 41766 45332 41804
rect 45612 41188 45668 41198
rect 45724 41188 45780 42478
rect 45612 41186 45780 41188
rect 45612 41134 45614 41186
rect 45666 41134 45780 41186
rect 45612 41132 45780 41134
rect 45612 41122 45668 41132
rect 45164 39566 45166 39618
rect 45218 39566 45220 39618
rect 45164 39554 45220 39566
rect 45276 41074 45332 41086
rect 45276 41022 45278 41074
rect 45330 41022 45332 41074
rect 45276 39396 45332 41022
rect 45836 41076 45892 41086
rect 45836 40982 45892 41020
rect 45724 40964 45780 40974
rect 45724 40870 45780 40908
rect 46172 40740 46228 47180
rect 47180 46674 47236 48076
rect 48188 48130 48244 48748
rect 48188 48078 48190 48130
rect 48242 48078 48244 48130
rect 48188 48020 48244 48078
rect 48188 47348 48244 47964
rect 47180 46622 47182 46674
rect 47234 46622 47236 46674
rect 46508 46564 46564 46574
rect 46508 46470 46564 46508
rect 47180 46564 47236 46622
rect 47964 47292 48244 47348
rect 48300 48802 48356 48814
rect 48300 48750 48302 48802
rect 48354 48750 48356 48802
rect 47740 46564 47796 46574
rect 47180 46562 47796 46564
rect 47180 46510 47742 46562
rect 47794 46510 47796 46562
rect 47180 46508 47796 46510
rect 46620 45332 46676 45342
rect 46620 44994 46676 45276
rect 46620 44942 46622 44994
rect 46674 44942 46676 44994
rect 46620 44930 46676 44942
rect 47068 44996 47124 45006
rect 47180 44996 47236 46508
rect 47740 46498 47796 46508
rect 47852 45108 47908 45118
rect 47964 45108 48020 47292
rect 48188 46676 48244 46686
rect 48188 46582 48244 46620
rect 48188 45220 48244 45230
rect 48300 45220 48356 48750
rect 48748 48356 48804 48366
rect 48860 48356 48916 48860
rect 48972 48850 49028 48860
rect 48748 48354 48916 48356
rect 48748 48302 48750 48354
rect 48802 48302 48916 48354
rect 48748 48300 48916 48302
rect 48748 48290 48804 48300
rect 49196 48244 49252 48972
rect 48860 48188 49252 48244
rect 49308 48244 49364 48254
rect 48748 47348 48804 47358
rect 48748 46900 48804 47292
rect 48636 46844 48804 46900
rect 48860 47234 48916 48188
rect 49308 48130 49364 48188
rect 49308 48078 49310 48130
rect 49362 48078 49364 48130
rect 49308 48066 49364 48078
rect 48972 48020 49028 48030
rect 48972 47926 49028 47964
rect 49644 47796 49700 49196
rect 48860 47182 48862 47234
rect 48914 47182 48916 47234
rect 48860 46900 48916 47182
rect 48636 46452 48692 46844
rect 48860 46834 48916 46844
rect 48972 47740 49700 47796
rect 49756 49026 49812 49038
rect 49756 48974 49758 49026
rect 49810 48974 49812 49026
rect 48748 46676 48804 46686
rect 48748 46582 48804 46620
rect 48636 46396 48804 46452
rect 48188 45218 48356 45220
rect 48188 45166 48190 45218
rect 48242 45166 48356 45218
rect 48188 45164 48356 45166
rect 48188 45154 48244 45164
rect 47852 45106 48020 45108
rect 47852 45054 47854 45106
rect 47906 45054 48020 45106
rect 47852 45052 48020 45054
rect 48300 45108 48356 45164
rect 48748 45220 48804 46396
rect 48972 45332 49028 47740
rect 49644 47570 49700 47582
rect 49644 47518 49646 47570
rect 49698 47518 49700 47570
rect 49084 47236 49140 47246
rect 49644 47236 49700 47518
rect 49084 47234 49700 47236
rect 49084 47182 49086 47234
rect 49138 47182 49700 47234
rect 49084 47180 49700 47182
rect 49084 47170 49140 47180
rect 49308 46564 49364 46574
rect 49308 45892 49364 46508
rect 49308 45826 49364 45836
rect 48748 45154 48804 45164
rect 48860 45276 49028 45332
rect 49084 45778 49140 45790
rect 49756 45780 49812 48974
rect 49980 49028 50036 49038
rect 49980 48466 50036 48972
rect 49980 48414 49982 48466
rect 50034 48414 50036 48466
rect 49980 48402 50036 48414
rect 49868 48242 49924 48254
rect 49868 48190 49870 48242
rect 49922 48190 49924 48242
rect 49868 47348 49924 48190
rect 49980 48244 50036 48254
rect 49980 47458 50036 48188
rect 49980 47406 49982 47458
rect 50034 47406 50036 47458
rect 49980 47394 50036 47406
rect 49868 47282 49924 47292
rect 49980 46564 50036 46574
rect 50092 46564 50148 49644
rect 50204 49252 50260 49262
rect 50204 48466 50260 49196
rect 50428 49252 50484 49262
rect 50540 49252 50596 49980
rect 51100 49924 51156 49934
rect 51324 49924 51380 51214
rect 51436 51268 51492 51326
rect 51660 51378 51716 51886
rect 51660 51326 51662 51378
rect 51714 51326 51716 51378
rect 51660 51314 51716 51326
rect 51436 51202 51492 51212
rect 51660 50596 51716 50606
rect 51100 49922 51380 49924
rect 51100 49870 51102 49922
rect 51154 49870 51380 49922
rect 51100 49868 51380 49870
rect 51436 50594 51716 50596
rect 51436 50542 51662 50594
rect 51714 50542 51716 50594
rect 51436 50540 51716 50542
rect 51100 49858 51156 49868
rect 50484 49196 50596 49252
rect 50428 49186 50484 49196
rect 50556 48636 50820 48646
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50556 48570 50820 48580
rect 50204 48414 50206 48466
rect 50258 48414 50260 48466
rect 50204 48402 50260 48414
rect 51100 48244 51156 48254
rect 51100 48242 51268 48244
rect 51100 48190 51102 48242
rect 51154 48190 51268 48242
rect 51100 48188 51268 48190
rect 51100 48178 51156 48188
rect 51212 47684 51268 48188
rect 51324 47684 51380 47694
rect 51212 47682 51380 47684
rect 51212 47630 51326 47682
rect 51378 47630 51380 47682
rect 51212 47628 51380 47630
rect 51324 47618 51380 47628
rect 51100 47570 51156 47582
rect 51100 47518 51102 47570
rect 51154 47518 51156 47570
rect 50428 47348 50484 47358
rect 50764 47348 50820 47358
rect 50428 47346 50820 47348
rect 50428 47294 50430 47346
rect 50482 47294 50766 47346
rect 50818 47294 50820 47346
rect 50428 47292 50820 47294
rect 50428 47282 50484 47292
rect 50764 47282 50820 47292
rect 50988 47234 51044 47246
rect 50988 47182 50990 47234
rect 51042 47182 51044 47234
rect 50556 47068 50820 47078
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50556 47002 50820 47012
rect 50316 46674 50372 46686
rect 50316 46622 50318 46674
rect 50370 46622 50372 46674
rect 50316 46564 50372 46622
rect 50988 46676 51044 47182
rect 51100 46786 51156 47518
rect 51436 47124 51492 50540
rect 51660 50530 51716 50540
rect 53228 49698 53284 49710
rect 53228 49646 53230 49698
rect 53282 49646 53284 49698
rect 51884 49138 51940 49150
rect 51884 49086 51886 49138
rect 51938 49086 51940 49138
rect 51884 48916 51940 49086
rect 53228 49140 53284 49646
rect 53228 49074 53284 49084
rect 51884 48850 51940 48860
rect 53004 48018 53060 48030
rect 53004 47966 53006 48018
rect 53058 47966 53060 48018
rect 51100 46734 51102 46786
rect 51154 46734 51156 46786
rect 51100 46722 51156 46734
rect 51212 47068 51492 47124
rect 51548 47682 51604 47694
rect 51548 47630 51550 47682
rect 51602 47630 51604 47682
rect 50988 46610 51044 46620
rect 49980 46562 50372 46564
rect 49980 46510 49982 46562
rect 50034 46510 50372 46562
rect 49980 46508 50372 46510
rect 49980 46498 50036 46508
rect 49084 45726 49086 45778
rect 49138 45726 49140 45778
rect 47068 44994 47236 44996
rect 47068 44942 47070 44994
rect 47122 44942 47236 44994
rect 47068 44940 47236 44942
rect 47516 44996 47572 45006
rect 47852 44996 47908 45052
rect 48300 45042 48356 45052
rect 47516 44994 47908 44996
rect 47516 44942 47518 44994
rect 47570 44942 47908 44994
rect 47516 44940 47908 44942
rect 48076 44994 48132 45006
rect 48076 44942 48078 44994
rect 48130 44942 48132 44994
rect 47068 43764 47124 44940
rect 46956 43708 47124 43764
rect 46284 43540 46340 43550
rect 46284 43538 46900 43540
rect 46284 43486 46286 43538
rect 46338 43486 46900 43538
rect 46284 43484 46900 43486
rect 46284 43474 46340 43484
rect 46844 41076 46900 43484
rect 46956 42756 47012 43708
rect 47516 43540 47572 44940
rect 48076 44660 48132 44942
rect 48748 44994 48804 45006
rect 48748 44942 48750 44994
rect 48802 44942 48804 44994
rect 48076 44604 48580 44660
rect 48524 44434 48580 44604
rect 48524 44382 48526 44434
rect 48578 44382 48580 44434
rect 48524 44370 48580 44382
rect 47516 43474 47572 43484
rect 46956 41972 47012 42700
rect 46956 41906 47012 41916
rect 47180 43428 47236 43438
rect 46844 41020 47012 41076
rect 45500 40684 46228 40740
rect 45388 39506 45444 39518
rect 45388 39454 45390 39506
rect 45442 39454 45444 39506
rect 45388 39396 45444 39454
rect 45332 39340 45444 39396
rect 45276 39330 45332 39340
rect 45276 36484 45332 36494
rect 45276 35700 45332 36428
rect 45276 35698 45444 35700
rect 45276 35646 45278 35698
rect 45330 35646 45444 35698
rect 45276 35644 45444 35646
rect 45276 35634 45332 35644
rect 44940 34802 45108 34804
rect 44940 34750 44942 34802
rect 44994 34750 45108 34802
rect 44940 34748 45108 34750
rect 44940 34738 44996 34748
rect 43820 34524 44100 34580
rect 45164 34690 45220 34702
rect 45164 34638 45166 34690
rect 45218 34638 45220 34690
rect 43820 34354 43876 34524
rect 43820 34302 43822 34354
rect 43874 34302 43876 34354
rect 43820 34290 43876 34302
rect 43708 34132 43764 34142
rect 43708 34038 43764 34076
rect 43820 33908 43876 33918
rect 43708 33906 43876 33908
rect 43708 33854 43822 33906
rect 43874 33854 43876 33906
rect 43708 33852 43876 33854
rect 43372 32786 43540 32788
rect 43372 32734 43374 32786
rect 43426 32734 43540 32786
rect 43372 32732 43540 32734
rect 43596 32788 43652 32798
rect 43372 32722 43428 32732
rect 43596 32694 43652 32732
rect 42924 32562 42980 32574
rect 42924 32510 42926 32562
rect 42978 32510 42980 32562
rect 42588 32450 42644 32462
rect 42588 32398 42590 32450
rect 42642 32398 42644 32450
rect 42588 32340 42644 32398
rect 42588 32274 42644 32284
rect 42924 32228 42980 32510
rect 43148 32562 43204 32574
rect 43596 32564 43652 32574
rect 43148 32510 43150 32562
rect 43202 32510 43204 32562
rect 43148 32340 43204 32510
rect 43148 32274 43204 32284
rect 43372 32562 43652 32564
rect 43372 32510 43598 32562
rect 43650 32510 43652 32562
rect 43372 32508 43652 32510
rect 42924 32162 42980 32172
rect 42812 31780 42868 31790
rect 42364 31724 42532 31780
rect 42252 31668 42308 31678
rect 42308 31612 42420 31668
rect 42252 31602 42308 31612
rect 42364 31554 42420 31612
rect 42364 31502 42366 31554
rect 42418 31502 42420 31554
rect 42364 31490 42420 31502
rect 42084 29708 42196 29764
rect 42028 29698 42084 29708
rect 41300 29484 41412 29540
rect 41692 29538 41860 29540
rect 41692 29486 41806 29538
rect 41858 29486 41860 29538
rect 41692 29484 41860 29486
rect 41244 29446 41300 29484
rect 41020 28866 41076 28878
rect 41020 28814 41022 28866
rect 41074 28814 41076 28866
rect 41020 28754 41076 28814
rect 41020 28702 41022 28754
rect 41074 28702 41076 28754
rect 41020 28690 41076 28702
rect 41132 28756 41188 28766
rect 41132 26514 41188 28700
rect 41356 28084 41412 28094
rect 41356 27300 41412 28028
rect 41356 27234 41412 27244
rect 41468 27076 41524 27114
rect 41468 27010 41524 27020
rect 41692 26908 41748 29484
rect 41804 29474 41860 29484
rect 42140 29540 42196 29550
rect 42140 29446 42196 29484
rect 41916 28756 41972 28766
rect 41916 28642 41972 28700
rect 41916 28590 41918 28642
rect 41970 28590 41972 28642
rect 41916 28578 41972 28590
rect 42476 28642 42532 31724
rect 42812 31686 42868 31724
rect 43372 31780 43428 32508
rect 43596 32498 43652 32508
rect 43708 32340 43764 33852
rect 43820 33842 43876 33852
rect 43372 31714 43428 31724
rect 43484 32284 43764 32340
rect 43932 33012 43988 33022
rect 43484 31778 43540 32284
rect 43484 31726 43486 31778
rect 43538 31726 43540 31778
rect 43484 31714 43540 31726
rect 43596 32116 43652 32126
rect 42700 31668 42756 31678
rect 42700 31574 42756 31612
rect 42812 31444 42868 31454
rect 42812 31220 42868 31388
rect 43372 31444 43428 31454
rect 43260 31220 43316 31230
rect 42812 31218 43316 31220
rect 42812 31166 42814 31218
rect 42866 31166 43262 31218
rect 43314 31166 43316 31218
rect 42812 31164 43316 31166
rect 42812 31154 42868 31164
rect 43260 31154 43316 31164
rect 43036 30996 43092 31006
rect 43036 30902 43092 30940
rect 42588 30212 42644 30222
rect 42588 30118 42644 30156
rect 42588 29764 42644 29774
rect 42588 29314 42644 29708
rect 42588 29262 42590 29314
rect 42642 29262 42644 29314
rect 42588 29250 42644 29262
rect 42924 28868 42980 28906
rect 42924 28802 42980 28812
rect 43372 28756 43428 31388
rect 43484 31220 43540 31230
rect 43596 31220 43652 32060
rect 43484 31218 43652 31220
rect 43484 31166 43486 31218
rect 43538 31166 43652 31218
rect 43484 31164 43652 31166
rect 43708 31780 43764 31790
rect 43484 31154 43540 31164
rect 43708 31108 43764 31724
rect 43820 31778 43876 31790
rect 43820 31726 43822 31778
rect 43874 31726 43876 31778
rect 43820 31444 43876 31726
rect 43820 31378 43876 31388
rect 43820 31220 43876 31230
rect 43820 31126 43876 31164
rect 43708 31014 43764 31052
rect 43260 28700 43428 28756
rect 43484 28756 43540 28766
rect 42476 28590 42478 28642
rect 42530 28590 42532 28642
rect 42476 28578 42532 28590
rect 42924 28644 42980 28654
rect 42924 28550 42980 28588
rect 41804 28530 41860 28542
rect 41804 28478 41806 28530
rect 41858 28478 41860 28530
rect 41804 28084 41860 28478
rect 43260 28420 43316 28700
rect 43484 28662 43540 28700
rect 43260 28354 43316 28364
rect 43372 28532 43428 28542
rect 41804 28018 41860 28028
rect 43372 28082 43428 28476
rect 43932 28420 43988 32956
rect 45164 32116 45220 34638
rect 45388 34130 45444 35644
rect 45500 34356 45556 40684
rect 46844 40290 46900 40302
rect 46844 40238 46846 40290
rect 46898 40238 46900 40290
rect 46172 39788 46788 39844
rect 45612 39620 45668 39630
rect 45612 38668 45668 39564
rect 46060 39508 46116 39518
rect 46060 39414 46116 39452
rect 46172 39394 46228 39788
rect 46732 39730 46788 39788
rect 46732 39678 46734 39730
rect 46786 39678 46788 39730
rect 46732 39666 46788 39678
rect 46172 39342 46174 39394
rect 46226 39342 46228 39394
rect 46172 39284 46228 39342
rect 46060 39228 46228 39284
rect 46284 39620 46340 39630
rect 45724 38836 45780 38874
rect 45724 38770 45780 38780
rect 45612 38612 46004 38668
rect 45948 38162 46004 38612
rect 45948 38110 45950 38162
rect 46002 38110 46004 38162
rect 45948 38098 46004 38110
rect 46060 36372 46116 39228
rect 46284 38836 46340 39564
rect 46844 39620 46900 40238
rect 46956 39620 47012 41020
rect 46956 39564 47124 39620
rect 46844 39554 46900 39564
rect 46396 39396 46452 39406
rect 46396 39394 46676 39396
rect 46396 39342 46398 39394
rect 46450 39342 46676 39394
rect 46396 39340 46676 39342
rect 46396 39330 46452 39340
rect 46396 39060 46452 39070
rect 46396 38966 46452 39004
rect 46284 38668 46340 38780
rect 46620 38834 46676 39340
rect 46956 39172 47012 39182
rect 46956 39058 47012 39116
rect 46956 39006 46958 39058
rect 47010 39006 47012 39058
rect 46956 38994 47012 39006
rect 47068 38946 47124 39564
rect 47068 38894 47070 38946
rect 47122 38894 47124 38946
rect 47068 38882 47124 38894
rect 46620 38782 46622 38834
rect 46674 38782 46676 38834
rect 46620 38770 46676 38782
rect 46172 38612 46340 38668
rect 47180 38668 47236 43372
rect 48300 43428 48356 43438
rect 48300 43334 48356 43372
rect 48748 42980 48804 44942
rect 48748 42914 48804 42924
rect 48860 42756 48916 45276
rect 48972 45108 49028 45118
rect 49084 45108 49140 45726
rect 49644 45724 49812 45780
rect 50204 45892 50260 45902
rect 49196 45668 49252 45678
rect 49196 45574 49252 45612
rect 49196 45108 49252 45118
rect 49084 45106 49252 45108
rect 49084 45054 49198 45106
rect 49250 45054 49252 45106
rect 49084 45052 49252 45054
rect 48972 45014 49028 45052
rect 49084 44660 49140 44670
rect 48972 44604 49084 44660
rect 48972 44322 49028 44604
rect 49084 44594 49140 44604
rect 48972 44270 48974 44322
rect 49026 44270 49028 44322
rect 48972 44258 49028 44270
rect 49084 43538 49140 43550
rect 49084 43486 49086 43538
rect 49138 43486 49140 43538
rect 48972 43428 49028 43438
rect 49084 43428 49140 43486
rect 49028 43372 49140 43428
rect 49196 43428 49252 45052
rect 49644 44436 49700 45724
rect 49868 45668 49924 45678
rect 49924 45612 50036 45668
rect 49868 45602 49924 45612
rect 49980 45330 50036 45612
rect 49980 45278 49982 45330
rect 50034 45278 50036 45330
rect 49980 45266 50036 45278
rect 50092 45220 50148 45230
rect 50092 45126 50148 45164
rect 49756 45106 49812 45118
rect 49756 45054 49758 45106
rect 49810 45054 49812 45106
rect 49756 44660 49812 45054
rect 49756 44594 49812 44604
rect 49644 44380 49812 44436
rect 49420 44210 49476 44222
rect 49420 44158 49422 44210
rect 49474 44158 49476 44210
rect 49308 43540 49364 43550
rect 49420 43540 49476 44158
rect 49644 44212 49700 44222
rect 49644 43650 49700 44156
rect 49644 43598 49646 43650
rect 49698 43598 49700 43650
rect 49644 43586 49700 43598
rect 49308 43538 49476 43540
rect 49308 43486 49310 43538
rect 49362 43486 49476 43538
rect 49308 43484 49476 43486
rect 49308 43474 49364 43484
rect 48972 43362 49028 43372
rect 49196 43362 49252 43372
rect 48748 42700 48916 42756
rect 48076 41972 48132 41982
rect 48076 41878 48132 41916
rect 47404 41858 47460 41870
rect 47404 41806 47406 41858
rect 47458 41806 47460 41858
rect 47404 40964 47460 41806
rect 48524 41188 48580 41198
rect 48412 41186 48580 41188
rect 48412 41134 48526 41186
rect 48578 41134 48580 41186
rect 48412 41132 48580 41134
rect 48412 40964 48468 41132
rect 48524 41122 48580 41132
rect 47404 40898 47460 40908
rect 48300 40962 48468 40964
rect 48300 40910 48414 40962
rect 48466 40910 48468 40962
rect 48300 40908 48468 40910
rect 47292 39060 47348 39070
rect 47292 38946 47348 39004
rect 47292 38894 47294 38946
rect 47346 38894 47348 38946
rect 47292 38882 47348 38894
rect 47180 38612 47348 38668
rect 46172 36484 46228 38612
rect 46172 36390 46228 36428
rect 46956 37156 47012 37166
rect 46844 36372 46900 36382
rect 46060 36306 46116 36316
rect 46284 36370 46900 36372
rect 46284 36318 46846 36370
rect 46898 36318 46900 36370
rect 46284 36316 46900 36318
rect 46284 35922 46340 36316
rect 46844 36306 46900 36316
rect 46284 35870 46286 35922
rect 46338 35870 46340 35922
rect 46284 35858 46340 35870
rect 46620 35812 46676 35822
rect 46956 35812 47012 37100
rect 46620 35810 47012 35812
rect 46620 35758 46622 35810
rect 46674 35758 47012 35810
rect 46620 35756 47012 35758
rect 46620 35746 46676 35756
rect 45948 35698 46004 35710
rect 45948 35646 45950 35698
rect 46002 35646 46004 35698
rect 45948 35364 46004 35646
rect 46284 35700 46340 35710
rect 46284 35606 46340 35644
rect 45948 35298 46004 35308
rect 45500 34290 45556 34300
rect 45388 34078 45390 34130
rect 45442 34078 45444 34130
rect 45388 34066 45444 34078
rect 46060 34020 46116 34030
rect 45500 34018 46116 34020
rect 45500 33966 46062 34018
rect 46114 33966 46116 34018
rect 45500 33964 46116 33966
rect 45500 33458 45556 33964
rect 46060 33954 46116 33964
rect 45500 33406 45502 33458
rect 45554 33406 45556 33458
rect 45500 33394 45556 33406
rect 45948 33684 46004 33694
rect 45612 33348 45668 33358
rect 45612 33254 45668 33292
rect 45948 33346 46004 33628
rect 45948 33294 45950 33346
rect 46002 33294 46004 33346
rect 45948 33282 46004 33294
rect 45164 32050 45220 32060
rect 45388 33234 45444 33246
rect 45388 33182 45390 33234
rect 45442 33182 45444 33234
rect 44156 31780 44212 31790
rect 44156 31686 44212 31724
rect 44940 31778 44996 31790
rect 44940 31726 44942 31778
rect 44994 31726 44996 31778
rect 44380 31556 44436 31566
rect 44380 31220 44436 31500
rect 44156 31218 44436 31220
rect 44156 31166 44382 31218
rect 44434 31166 44436 31218
rect 44156 31164 44436 31166
rect 44044 31108 44100 31118
rect 44044 31014 44100 31052
rect 44044 28644 44100 28654
rect 44156 28644 44212 31164
rect 44380 31154 44436 31164
rect 44828 31108 44884 31118
rect 44828 31014 44884 31052
rect 44716 30994 44772 31006
rect 44716 30942 44718 30994
rect 44770 30942 44772 30994
rect 44044 28642 44212 28644
rect 44044 28590 44046 28642
rect 44098 28590 44212 28642
rect 44044 28588 44212 28590
rect 44268 29426 44324 29438
rect 44268 29374 44270 29426
rect 44322 29374 44324 29426
rect 44268 28644 44324 29374
rect 44604 28644 44660 28654
rect 44268 28588 44604 28644
rect 44044 28578 44100 28588
rect 44604 28578 44660 28588
rect 43932 28364 44324 28420
rect 43372 28030 43374 28082
rect 43426 28030 43428 28082
rect 43372 28018 43428 28030
rect 43708 27748 43764 27758
rect 43708 27654 43764 27692
rect 43932 27746 43988 27758
rect 43932 27694 43934 27746
rect 43986 27694 43988 27746
rect 43932 27636 43988 27694
rect 44156 27636 44212 27646
rect 43932 27634 44212 27636
rect 43932 27582 44158 27634
rect 44210 27582 44212 27634
rect 43932 27580 44212 27582
rect 44156 27570 44212 27580
rect 42476 27244 43204 27300
rect 41132 26462 41134 26514
rect 41186 26462 41188 26514
rect 41132 26450 41188 26462
rect 41468 26852 41748 26908
rect 42028 27186 42084 27198
rect 42028 27134 42030 27186
rect 42082 27134 42084 27186
rect 42028 26964 42084 27134
rect 41020 26402 41076 26414
rect 41020 26350 41022 26402
rect 41074 26350 41076 26402
rect 41020 26292 41076 26350
rect 41020 26236 41412 26292
rect 41356 26180 41412 26236
rect 40908 26124 41188 26180
rect 40796 25564 41076 25620
rect 40796 25396 40852 25406
rect 40796 24050 40852 25340
rect 40796 23998 40798 24050
rect 40850 23998 40852 24050
rect 40796 23986 40852 23998
rect 40908 21924 40964 21934
rect 40908 21586 40964 21868
rect 40908 21534 40910 21586
rect 40962 21534 40964 21586
rect 40908 21522 40964 21534
rect 41020 21140 41076 25564
rect 41132 25506 41188 26124
rect 41132 25454 41134 25506
rect 41186 25454 41188 25506
rect 41132 25442 41188 25454
rect 41244 26066 41300 26078
rect 41244 26014 41246 26066
rect 41298 26014 41300 26066
rect 41244 24612 41300 26014
rect 41244 24546 41300 24556
rect 41356 23938 41412 26124
rect 41356 23886 41358 23938
rect 41410 23886 41412 23938
rect 41356 22820 41412 23886
rect 41356 22754 41412 22764
rect 41244 22372 41300 22382
rect 41244 22278 41300 22316
rect 41468 22260 41524 26852
rect 42028 25620 42084 26908
rect 42140 27074 42196 27086
rect 42140 27022 42142 27074
rect 42194 27022 42196 27074
rect 42140 26180 42196 27022
rect 42476 27074 42532 27244
rect 42476 27022 42478 27074
rect 42530 27022 42532 27074
rect 42476 27010 42532 27022
rect 43036 27076 43092 27086
rect 42364 26516 42420 26526
rect 42364 26422 42420 26460
rect 42140 26114 42196 26124
rect 42924 26180 42980 26190
rect 42924 26086 42980 26124
rect 42588 25620 42644 25630
rect 42028 25618 42644 25620
rect 42028 25566 42030 25618
rect 42082 25566 42590 25618
rect 42642 25566 42644 25618
rect 42028 25564 42644 25566
rect 42028 25554 42084 25564
rect 42588 25554 42644 25564
rect 41580 25506 41636 25518
rect 41580 25454 41582 25506
rect 41634 25454 41636 25506
rect 41580 25284 41636 25454
rect 43036 25506 43092 27020
rect 43036 25454 43038 25506
rect 43090 25454 43092 25506
rect 42252 25284 42308 25294
rect 41580 25228 42084 25284
rect 42028 24724 42084 25228
rect 42252 25190 42308 25228
rect 42252 24724 42308 24734
rect 42028 24668 42252 24724
rect 41692 23268 41748 23278
rect 42028 23268 42084 24668
rect 42252 24630 42308 24668
rect 42140 24500 42196 24510
rect 42196 24444 42308 24500
rect 42140 24434 42196 24444
rect 41692 23266 42084 23268
rect 41692 23214 41694 23266
rect 41746 23214 42030 23266
rect 42082 23214 42084 23266
rect 41692 23212 42084 23214
rect 41692 23202 41748 23212
rect 42028 23202 42084 23212
rect 42140 23044 42196 23054
rect 42140 22950 42196 22988
rect 41468 22194 41524 22204
rect 41692 22370 41748 22382
rect 41692 22318 41694 22370
rect 41746 22318 41748 22370
rect 41692 22148 41748 22318
rect 41692 22082 41748 22092
rect 41356 21924 41412 21934
rect 41412 21868 41748 21924
rect 41356 21858 41412 21868
rect 41692 21810 41748 21868
rect 41692 21758 41694 21810
rect 41746 21758 41748 21810
rect 41692 21746 41748 21758
rect 41580 21700 41636 21710
rect 41132 21588 41188 21598
rect 41132 21494 41188 21532
rect 41244 21364 41300 21374
rect 41244 21270 41300 21308
rect 41076 21084 41412 21140
rect 41020 21074 41076 21084
rect 41020 20914 41076 20926
rect 41020 20862 41022 20914
rect 41074 20862 41076 20914
rect 40908 19908 40964 19918
rect 40908 19814 40964 19852
rect 41020 18452 41076 20862
rect 41356 20020 41412 21084
rect 41580 20802 41636 21644
rect 41580 20750 41582 20802
rect 41634 20750 41636 20802
rect 41580 20738 41636 20750
rect 42140 21476 42196 21486
rect 42252 21476 42308 24444
rect 42588 23826 42644 23838
rect 42588 23774 42590 23826
rect 42642 23774 42644 23826
rect 42588 23492 42644 23774
rect 42588 23426 42644 23436
rect 42812 23154 42868 23166
rect 42812 23102 42814 23154
rect 42866 23102 42868 23154
rect 42700 23044 42756 23054
rect 42812 23044 42868 23102
rect 43036 23154 43092 25454
rect 43148 26964 43204 27244
rect 44268 27298 44324 28364
rect 44492 27746 44548 27758
rect 44492 27694 44494 27746
rect 44546 27694 44548 27746
rect 44492 27636 44548 27694
rect 44268 27246 44270 27298
rect 44322 27246 44324 27298
rect 44268 27234 44324 27246
rect 44380 27634 44548 27636
rect 44380 27582 44494 27634
rect 44546 27582 44548 27634
rect 44380 27580 44548 27582
rect 43708 27074 43764 27086
rect 43708 27022 43710 27074
rect 43762 27022 43764 27074
rect 43372 26964 43428 26974
rect 43148 26962 43428 26964
rect 43148 26910 43374 26962
rect 43426 26910 43428 26962
rect 43148 26908 43428 26910
rect 43148 25506 43204 26908
rect 43372 26898 43428 26908
rect 43708 26964 43764 27022
rect 43708 26402 43764 26908
rect 43708 26350 43710 26402
rect 43762 26350 43764 26402
rect 43708 26338 43764 26350
rect 43932 27074 43988 27086
rect 43932 27022 43934 27074
rect 43986 27022 43988 27074
rect 43148 25454 43150 25506
rect 43202 25454 43204 25506
rect 43148 25060 43204 25454
rect 43148 24994 43204 25004
rect 43260 26290 43316 26302
rect 43260 26238 43262 26290
rect 43314 26238 43316 26290
rect 43260 26180 43316 26238
rect 43932 26180 43988 27022
rect 44156 27076 44212 27086
rect 44156 26982 44212 27020
rect 43260 26124 43988 26180
rect 43260 24834 43316 26124
rect 43260 24782 43262 24834
rect 43314 24782 43316 24834
rect 43036 23102 43038 23154
rect 43090 23102 43092 23154
rect 42924 23044 42980 23054
rect 42812 22988 42924 23044
rect 42588 22932 42644 22942
rect 42588 22838 42644 22876
rect 42700 22596 42756 22988
rect 42924 22978 42980 22988
rect 42812 22596 42868 22606
rect 42700 22594 42868 22596
rect 42700 22542 42814 22594
rect 42866 22542 42868 22594
rect 42700 22540 42868 22542
rect 42812 22530 42868 22540
rect 42476 22370 42532 22382
rect 42476 22318 42478 22370
rect 42530 22318 42532 22370
rect 42364 22258 42420 22270
rect 42364 22206 42366 22258
rect 42418 22206 42420 22258
rect 42364 22148 42420 22206
rect 42476 22148 42532 22318
rect 42700 22372 42756 22382
rect 42700 22278 42756 22316
rect 42700 22148 42756 22158
rect 42476 22092 42700 22148
rect 42364 22082 42420 22092
rect 42700 22082 42756 22092
rect 42140 21474 42308 21476
rect 42140 21422 42142 21474
rect 42194 21422 42308 21474
rect 42140 21420 42308 21422
rect 42812 21812 42868 21822
rect 41356 20018 41748 20020
rect 41356 19966 41358 20018
rect 41410 19966 41748 20018
rect 41356 19964 41748 19966
rect 41356 19954 41412 19964
rect 41692 19346 41748 19964
rect 41692 19294 41694 19346
rect 41746 19294 41748 19346
rect 41692 19282 41748 19294
rect 42140 19010 42196 21420
rect 42812 21364 42868 21756
rect 43036 21700 43092 23102
rect 43036 21634 43092 21644
rect 43148 24612 43204 24622
rect 43148 23938 43204 24556
rect 43148 23886 43150 23938
rect 43202 23886 43204 23938
rect 42812 21028 42868 21308
rect 42700 21026 42868 21028
rect 42700 20974 42814 21026
rect 42866 20974 42868 21026
rect 42700 20972 42868 20974
rect 42140 18958 42142 19010
rect 42194 18958 42196 19010
rect 42140 18900 42196 18958
rect 42140 18834 42196 18844
rect 42364 20578 42420 20590
rect 42364 20526 42366 20578
rect 42418 20526 42420 20578
rect 42028 18564 42084 18574
rect 42364 18564 42420 20526
rect 42700 20130 42756 20972
rect 42812 20962 42868 20972
rect 42700 20078 42702 20130
rect 42754 20078 42756 20130
rect 42700 20066 42756 20078
rect 43036 20804 43092 20814
rect 43148 20804 43204 23886
rect 43260 23380 43316 24782
rect 44044 25282 44100 25294
rect 44044 25230 44046 25282
rect 44098 25230 44100 25282
rect 44044 25060 44100 25230
rect 43484 24724 43540 24734
rect 43484 24612 43540 24668
rect 43932 24612 43988 24622
rect 43484 24610 43988 24612
rect 43484 24558 43934 24610
rect 43986 24558 43988 24610
rect 43484 24556 43988 24558
rect 43596 23828 43652 23838
rect 43596 23734 43652 23772
rect 43260 23314 43316 23324
rect 43484 23714 43540 23726
rect 43484 23662 43486 23714
rect 43538 23662 43540 23714
rect 43484 23156 43540 23662
rect 43260 22820 43316 22830
rect 43260 22482 43316 22764
rect 43260 22430 43262 22482
rect 43314 22430 43316 22482
rect 43260 22418 43316 22430
rect 43484 22372 43540 23100
rect 43484 22306 43540 22316
rect 43596 23492 43652 23502
rect 43596 21812 43652 23436
rect 43820 22148 43876 22158
rect 43820 22054 43876 22092
rect 43932 21924 43988 24556
rect 44044 23828 44100 25004
rect 44044 23734 44100 23772
rect 44156 23156 44212 23166
rect 44156 23062 44212 23100
rect 44268 22148 44324 22158
rect 44268 22054 44324 22092
rect 43596 21718 43652 21756
rect 43820 21868 43988 21924
rect 43484 21700 43540 21710
rect 43484 20916 43540 21644
rect 43820 21364 43876 21868
rect 44044 21698 44100 21710
rect 44044 21646 44046 21698
rect 44098 21646 44100 21698
rect 43932 21588 43988 21598
rect 43932 21494 43988 21532
rect 44044 21364 44100 21646
rect 44268 21364 44324 21374
rect 44380 21364 44436 27580
rect 44492 27570 44548 27580
rect 44716 26908 44772 30942
rect 44940 29876 44996 31726
rect 45164 31556 45220 31566
rect 45220 31500 45332 31556
rect 45164 31490 45220 31500
rect 45052 31108 45108 31118
rect 45052 31106 45220 31108
rect 45052 31054 45054 31106
rect 45106 31054 45220 31106
rect 45052 31052 45220 31054
rect 45052 31042 45108 31052
rect 45164 30996 45220 31052
rect 45164 30930 45220 30940
rect 45276 30100 45332 31500
rect 45164 30044 45332 30100
rect 44940 29820 45108 29876
rect 44940 29652 44996 29662
rect 44940 29538 44996 29596
rect 44940 29486 44942 29538
rect 44994 29486 44996 29538
rect 44940 29474 44996 29486
rect 44940 28642 44996 28654
rect 44940 28590 44942 28642
rect 44994 28590 44996 28642
rect 44940 28082 44996 28590
rect 44940 28030 44942 28082
rect 44994 28030 44996 28082
rect 44940 27634 44996 28030
rect 44940 27582 44942 27634
rect 44994 27582 44996 27634
rect 44940 27570 44996 27582
rect 45052 28644 45108 29820
rect 44604 26852 44772 26908
rect 44604 23604 44660 26852
rect 45052 26290 45108 28588
rect 45164 28530 45220 30044
rect 45164 28478 45166 28530
rect 45218 28478 45220 28530
rect 45164 28466 45220 28478
rect 45276 27748 45332 27758
rect 45276 26908 45332 27692
rect 45388 27524 45444 33182
rect 45612 32452 45668 32462
rect 45612 31890 45668 32396
rect 45612 31838 45614 31890
rect 45666 31838 45668 31890
rect 45612 31826 45668 31838
rect 47292 30212 47348 38612
rect 48188 37154 48244 37166
rect 48188 37102 48190 37154
rect 48242 37102 48244 37154
rect 48188 37044 48244 37102
rect 48188 36978 48244 36988
rect 47292 30146 47348 30156
rect 47404 34692 47460 34702
rect 47068 30100 47124 30110
rect 47068 29316 47124 30044
rect 46956 29314 47124 29316
rect 46956 29262 47070 29314
rect 47122 29262 47124 29314
rect 46956 29260 47124 29262
rect 46508 28756 46564 28766
rect 45500 27748 45556 27758
rect 45500 27654 45556 27692
rect 45388 27468 46452 27524
rect 45500 27188 45556 27198
rect 45276 26852 45444 26908
rect 45052 26238 45054 26290
rect 45106 26238 45108 26290
rect 45052 26226 45108 26238
rect 45388 23940 45444 26852
rect 45500 25620 45556 27132
rect 45836 26178 45892 26190
rect 45836 26126 45838 26178
rect 45890 26126 45892 26178
rect 45724 25732 45780 25742
rect 45836 25732 45892 26126
rect 45724 25730 45892 25732
rect 45724 25678 45726 25730
rect 45778 25678 45892 25730
rect 45724 25676 45892 25678
rect 45724 25666 45780 25676
rect 45500 25618 45668 25620
rect 45500 25566 45502 25618
rect 45554 25566 45668 25618
rect 45500 25564 45668 25566
rect 45500 25554 45556 25564
rect 45612 25508 45668 25564
rect 45836 25508 45892 25518
rect 45612 25506 45892 25508
rect 45612 25454 45838 25506
rect 45890 25454 45892 25506
rect 45612 25452 45892 25454
rect 45836 25442 45892 25452
rect 46060 25508 46116 25518
rect 45724 24722 45780 24734
rect 45724 24670 45726 24722
rect 45778 24670 45780 24722
rect 45724 24162 45780 24670
rect 45724 24110 45726 24162
rect 45778 24110 45780 24162
rect 45724 24098 45780 24110
rect 45388 23884 45556 23940
rect 44604 23538 44660 23548
rect 44828 23828 44884 23838
rect 44492 23044 44548 23054
rect 44492 22950 44548 22988
rect 43820 21308 43988 21364
rect 44044 21362 44436 21364
rect 44044 21310 44270 21362
rect 44322 21310 44436 21362
rect 44044 21308 44436 21310
rect 44492 22148 44548 22158
rect 44492 21474 44548 22092
rect 44492 21422 44494 21474
rect 44546 21422 44548 21474
rect 43484 20914 43876 20916
rect 43484 20862 43486 20914
rect 43538 20862 43876 20914
rect 43484 20860 43876 20862
rect 43484 20850 43540 20860
rect 43036 20802 43204 20804
rect 43036 20750 43038 20802
rect 43090 20750 43204 20802
rect 43036 20748 43204 20750
rect 43260 20802 43316 20814
rect 43260 20750 43262 20802
rect 43314 20750 43316 20802
rect 43036 20020 43092 20748
rect 43260 20244 43316 20750
rect 43820 20690 43876 20860
rect 43820 20638 43822 20690
rect 43874 20638 43876 20690
rect 43820 20626 43876 20638
rect 43932 20468 43988 21308
rect 44268 21298 44324 21308
rect 44492 20804 44548 21422
rect 44828 21140 44884 23772
rect 45388 23714 45444 23726
rect 45388 23662 45390 23714
rect 45442 23662 45444 23714
rect 45388 23492 45444 23662
rect 45388 23426 45444 23436
rect 45500 23268 45556 23884
rect 45612 23826 45668 23838
rect 45612 23774 45614 23826
rect 45666 23774 45668 23826
rect 45612 23380 45668 23774
rect 45724 23714 45780 23726
rect 45724 23662 45726 23714
rect 45778 23662 45780 23714
rect 45724 23604 45780 23662
rect 45724 23538 45780 23548
rect 46060 23548 46116 25452
rect 46284 25506 46340 25518
rect 46284 25454 46286 25506
rect 46338 25454 46340 25506
rect 46172 25396 46228 25406
rect 46172 24946 46228 25340
rect 46172 24894 46174 24946
rect 46226 24894 46228 24946
rect 46172 24882 46228 24894
rect 46284 24946 46340 25454
rect 46396 25172 46452 27468
rect 46396 25106 46452 25116
rect 46284 24894 46286 24946
rect 46338 24894 46340 24946
rect 46284 24882 46340 24894
rect 46396 24722 46452 24734
rect 46396 24670 46398 24722
rect 46450 24670 46452 24722
rect 46172 23940 46228 23950
rect 46172 23846 46228 23884
rect 46060 23492 46340 23548
rect 45612 23314 45668 23324
rect 45164 23212 45556 23268
rect 45052 22148 45108 22158
rect 45052 22054 45108 22092
rect 45164 21588 45220 23212
rect 45724 23154 45780 23166
rect 45724 23102 45726 23154
rect 45778 23102 45780 23154
rect 45276 23044 45332 23054
rect 45724 23044 45780 23102
rect 45276 23042 45780 23044
rect 45276 22990 45278 23042
rect 45330 22990 45780 23042
rect 45276 22988 45780 22990
rect 45276 22978 45332 22988
rect 45724 22370 45780 22988
rect 45724 22318 45726 22370
rect 45778 22318 45780 22370
rect 45388 22260 45444 22270
rect 45388 22166 45444 22204
rect 45388 21924 45444 21934
rect 45724 21924 45780 22318
rect 46284 22932 46340 23492
rect 46396 23380 46452 24670
rect 46396 23314 46452 23324
rect 46284 22260 46340 22876
rect 46284 22194 46340 22204
rect 45444 21868 45780 21924
rect 45388 21858 45444 21868
rect 45276 21588 45332 21598
rect 45164 21532 45276 21588
rect 44940 21474 44996 21486
rect 44940 21422 44942 21474
rect 44994 21422 44996 21474
rect 44940 21364 44996 21422
rect 45276 21476 45332 21532
rect 45388 21476 45444 21486
rect 45276 21474 45444 21476
rect 45276 21422 45390 21474
rect 45442 21422 45444 21474
rect 45276 21420 45444 21422
rect 44940 21362 45220 21364
rect 44940 21310 44942 21362
rect 44994 21310 45220 21362
rect 44940 21308 45220 21310
rect 44940 21270 44996 21308
rect 44828 21084 45108 21140
rect 44492 20748 44996 20804
rect 44940 20692 44996 20748
rect 44940 20598 44996 20636
rect 44156 20580 44212 20590
rect 44828 20580 44884 20590
rect 44156 20578 44884 20580
rect 44156 20526 44158 20578
rect 44210 20526 44830 20578
rect 44882 20526 44884 20578
rect 44156 20524 44884 20526
rect 44156 20514 44212 20524
rect 43260 20178 43316 20188
rect 43820 20412 43988 20468
rect 43708 20020 43764 20030
rect 43036 20018 43764 20020
rect 43036 19966 43710 20018
rect 43762 19966 43764 20018
rect 43036 19964 43764 19966
rect 43708 19954 43764 19964
rect 43372 18900 43428 18910
rect 42588 18564 42644 18574
rect 42084 18508 42196 18564
rect 42364 18508 42588 18564
rect 42028 18498 42084 18508
rect 41020 18386 41076 18396
rect 41804 18452 41860 18462
rect 41804 18358 41860 18396
rect 41916 18340 41972 18350
rect 40684 18172 41300 18228
rect 40460 17668 40516 17678
rect 40460 17574 40516 17612
rect 41244 17108 41300 18172
rect 41244 17106 41636 17108
rect 41244 17054 41246 17106
rect 41298 17054 41636 17106
rect 41244 17052 41636 17054
rect 41244 17042 41300 17052
rect 41580 16882 41636 17052
rect 41916 17106 41972 18284
rect 42140 17668 42196 18508
rect 42252 18452 42308 18462
rect 42252 18358 42308 18396
rect 42252 17668 42308 17678
rect 42140 17666 42308 17668
rect 42140 17614 42254 17666
rect 42306 17614 42308 17666
rect 42140 17612 42308 17614
rect 42252 17602 42308 17612
rect 41916 17054 41918 17106
rect 41970 17054 41972 17106
rect 41916 17042 41972 17054
rect 42028 17554 42084 17566
rect 42028 17502 42030 17554
rect 42082 17502 42084 17554
rect 42028 16996 42084 17502
rect 41580 16830 41582 16882
rect 41634 16830 41636 16882
rect 41580 16772 41636 16830
rect 41692 16828 41972 16884
rect 41692 16772 41748 16828
rect 41580 16716 41748 16772
rect 41804 16658 41860 16670
rect 41804 16606 41806 16658
rect 41858 16606 41860 16658
rect 40460 16210 40516 16222
rect 40460 16158 40462 16210
rect 40514 16158 40516 16210
rect 40460 15148 40516 16158
rect 41020 16212 41076 16222
rect 40796 16100 40852 16110
rect 40796 16006 40852 16044
rect 40684 15988 40740 15998
rect 40684 15894 40740 15932
rect 41020 15538 41076 16156
rect 41020 15486 41022 15538
rect 41074 15486 41076 15538
rect 40460 15092 40628 15148
rect 40908 15092 40964 15102
rect 40348 12338 40404 12348
rect 40460 13300 40516 13310
rect 39900 11676 40292 11732
rect 39900 10834 39956 11676
rect 40460 11618 40516 13244
rect 40572 12628 40628 15092
rect 40684 15090 40964 15092
rect 40684 15038 40910 15090
rect 40962 15038 40964 15090
rect 40684 15036 40964 15038
rect 40684 14644 40740 15036
rect 40908 15026 40964 15036
rect 40684 14530 40740 14588
rect 40684 14478 40686 14530
rect 40738 14478 40740 14530
rect 40684 14466 40740 14478
rect 41020 14530 41076 15486
rect 41468 15876 41524 15886
rect 41468 15426 41524 15820
rect 41468 15374 41470 15426
rect 41522 15374 41524 15426
rect 41468 15362 41524 15374
rect 41244 15316 41300 15354
rect 41244 15250 41300 15260
rect 41804 15148 41860 16606
rect 41132 15092 41860 15148
rect 41132 14642 41188 15092
rect 41916 14644 41972 16828
rect 42028 16882 42084 16940
rect 42028 16830 42030 16882
rect 42082 16830 42084 16882
rect 42028 16818 42084 16830
rect 42364 16882 42420 16894
rect 42364 16830 42366 16882
rect 42418 16830 42420 16882
rect 42364 16436 42420 16830
rect 42588 16660 42644 18508
rect 42924 18340 42980 18350
rect 42924 18246 42980 18284
rect 43260 18340 43316 18350
rect 43260 17668 43316 18284
rect 42812 17666 43316 17668
rect 42812 17614 43262 17666
rect 43314 17614 43316 17666
rect 42812 17612 43316 17614
rect 42700 16996 42756 17006
rect 42700 16902 42756 16940
rect 42812 16994 42868 17612
rect 43260 17602 43316 17612
rect 42812 16942 42814 16994
rect 42866 16942 42868 16994
rect 42812 16930 42868 16942
rect 42924 17442 42980 17454
rect 42924 17390 42926 17442
rect 42978 17390 42980 17442
rect 42588 16604 42756 16660
rect 42140 16380 42644 16436
rect 42140 15314 42196 16380
rect 42588 16098 42644 16380
rect 42588 16046 42590 16098
rect 42642 16046 42644 16098
rect 42588 16034 42644 16046
rect 42364 15428 42420 15438
rect 42364 15334 42420 15372
rect 42140 15262 42142 15314
rect 42194 15262 42196 15314
rect 42140 15250 42196 15262
rect 42252 15314 42308 15326
rect 42252 15262 42254 15314
rect 42306 15262 42308 15314
rect 42252 15148 42308 15262
rect 42476 15316 42532 15326
rect 42476 15222 42532 15260
rect 42588 15314 42644 15326
rect 42588 15262 42590 15314
rect 42642 15262 42644 15314
rect 41132 14590 41134 14642
rect 41186 14590 41188 14642
rect 41132 14578 41188 14590
rect 41804 14588 41972 14644
rect 42140 15092 42308 15148
rect 41020 14478 41022 14530
rect 41074 14478 41076 14530
rect 41020 14466 41076 14478
rect 41244 14530 41300 14542
rect 41244 14478 41246 14530
rect 41298 14478 41300 14530
rect 40796 14308 40852 14318
rect 40796 14214 40852 14252
rect 41244 14308 41300 14478
rect 41244 14242 41300 14252
rect 40572 12572 41524 12628
rect 41020 12404 41076 12414
rect 40460 11566 40462 11618
rect 40514 11566 40516 11618
rect 40460 11554 40516 11566
rect 40908 12348 41020 12404
rect 41076 12348 41300 12404
rect 39900 10782 39902 10834
rect 39954 10782 39956 10834
rect 39900 10386 39956 10782
rect 39900 10334 39902 10386
rect 39954 10334 39956 10386
rect 39900 10322 39956 10334
rect 40796 11396 40852 11406
rect 40796 11170 40852 11340
rect 40796 11118 40798 11170
rect 40850 11118 40852 11170
rect 39900 9716 39956 9726
rect 39900 9156 39956 9660
rect 40460 9714 40516 9726
rect 40460 9662 40462 9714
rect 40514 9662 40516 9714
rect 39900 9042 39956 9100
rect 39900 8990 39902 9042
rect 39954 8990 39956 9042
rect 39900 8978 39956 8990
rect 40124 9602 40180 9614
rect 40124 9550 40126 9602
rect 40178 9550 40180 9602
rect 40124 9044 40180 9550
rect 40124 8978 40180 8988
rect 40348 9044 40404 9054
rect 40460 9044 40516 9662
rect 40348 9042 40516 9044
rect 40348 8990 40350 9042
rect 40402 8990 40516 9042
rect 40348 8988 40516 8990
rect 40348 8484 40404 8988
rect 40348 8418 40404 8428
rect 40348 7474 40404 7486
rect 40348 7422 40350 7474
rect 40402 7422 40404 7474
rect 40348 7252 40404 7422
rect 40796 7476 40852 11118
rect 40796 7410 40852 7420
rect 40908 7700 40964 12348
rect 41020 12310 41076 12348
rect 41020 11618 41076 11630
rect 41020 11566 41022 11618
rect 41074 11566 41076 11618
rect 41020 10610 41076 11566
rect 41244 11506 41300 12348
rect 41244 11454 41246 11506
rect 41298 11454 41300 11506
rect 41244 11442 41300 11454
rect 41020 10558 41022 10610
rect 41074 10558 41076 10610
rect 41020 10052 41076 10558
rect 41020 9986 41076 9996
rect 41468 9828 41524 12572
rect 41580 12404 41636 12414
rect 41580 12178 41636 12348
rect 41580 12126 41582 12178
rect 41634 12126 41636 12178
rect 41580 12114 41636 12126
rect 41804 11396 41860 14588
rect 41916 14420 41972 14430
rect 41916 14326 41972 14364
rect 41916 14196 41972 14206
rect 42140 14196 42196 15092
rect 42588 14420 42644 15262
rect 42588 14354 42644 14364
rect 42252 14308 42308 14318
rect 42252 14214 42308 14252
rect 41972 14140 42196 14196
rect 41916 13186 41972 14140
rect 41916 13134 41918 13186
rect 41970 13134 41972 13186
rect 41916 13122 41972 13134
rect 42252 12964 42308 12974
rect 42028 12738 42084 12750
rect 42028 12686 42030 12738
rect 42082 12686 42084 12738
rect 42028 11618 42084 12686
rect 42028 11566 42030 11618
rect 42082 11566 42084 11618
rect 42028 11554 42084 11566
rect 41916 11396 41972 11406
rect 41804 11340 41916 11396
rect 41916 11302 41972 11340
rect 42252 11394 42308 12908
rect 42364 12066 42420 12078
rect 42364 12014 42366 12066
rect 42418 12014 42420 12066
rect 42364 11508 42420 12014
rect 42476 11508 42532 11518
rect 42364 11506 42532 11508
rect 42364 11454 42478 11506
rect 42530 11454 42532 11506
rect 42364 11452 42532 11454
rect 42476 11442 42532 11452
rect 42252 11342 42254 11394
rect 42306 11342 42308 11394
rect 42252 11330 42308 11342
rect 42588 11282 42644 11294
rect 42588 11230 42590 11282
rect 42642 11230 42644 11282
rect 41580 10498 41636 10510
rect 41580 10446 41582 10498
rect 41634 10446 41636 10498
rect 41580 10164 41636 10446
rect 42588 10388 42644 11230
rect 42700 10834 42756 16604
rect 42924 16212 42980 17390
rect 42924 16146 42980 16156
rect 43148 16212 43204 16222
rect 42924 15986 42980 15998
rect 42924 15934 42926 15986
rect 42978 15934 42980 15986
rect 42812 15874 42868 15886
rect 42812 15822 42814 15874
rect 42866 15822 42868 15874
rect 42812 15316 42868 15822
rect 42812 14420 42868 15260
rect 42924 15652 42980 15934
rect 42924 14644 42980 15596
rect 43148 15204 43204 16156
rect 43260 15764 43316 15774
rect 43260 15538 43316 15708
rect 43260 15486 43262 15538
rect 43314 15486 43316 15538
rect 43260 15474 43316 15486
rect 43372 15316 43428 18844
rect 43484 15652 43540 15662
rect 43484 15538 43540 15596
rect 43484 15486 43486 15538
rect 43538 15486 43540 15538
rect 43484 15474 43540 15486
rect 43148 15138 43204 15148
rect 43260 15260 43428 15316
rect 43708 15316 43764 15326
rect 42924 14588 43204 14644
rect 43036 14420 43092 14430
rect 42812 14418 43092 14420
rect 42812 14366 43038 14418
rect 43090 14366 43092 14418
rect 42812 14364 43092 14366
rect 43036 14354 43092 14364
rect 43148 12964 43204 14588
rect 43148 12898 43204 12908
rect 42700 10782 42702 10834
rect 42754 10782 42756 10834
rect 42700 10770 42756 10782
rect 43260 10724 43316 15260
rect 43708 15222 43764 15260
rect 43596 15202 43652 15214
rect 43596 15150 43598 15202
rect 43650 15150 43652 15202
rect 43596 15148 43652 15150
rect 43372 15092 43428 15102
rect 43596 15092 43764 15148
rect 43372 14530 43428 15036
rect 43708 15026 43764 15036
rect 43372 14478 43374 14530
rect 43426 14478 43428 14530
rect 43372 14466 43428 14478
rect 43708 12964 43764 12974
rect 43708 12850 43764 12908
rect 43708 12798 43710 12850
rect 43762 12798 43764 12850
rect 43708 12786 43764 12798
rect 43260 10668 43428 10724
rect 42812 10610 42868 10622
rect 42812 10558 42814 10610
rect 42866 10558 42868 10610
rect 42812 10500 42868 10558
rect 43260 10500 43316 10510
rect 42812 10498 43316 10500
rect 42812 10446 43262 10498
rect 43314 10446 43316 10498
rect 42812 10444 43316 10446
rect 42700 10388 42756 10398
rect 42588 10332 42700 10388
rect 42700 10294 42756 10332
rect 41692 10164 41748 10174
rect 41580 10108 41692 10164
rect 41020 9826 41524 9828
rect 41020 9774 41470 9826
rect 41522 9774 41524 9826
rect 41020 9772 41524 9774
rect 41020 8258 41076 9772
rect 41468 9762 41524 9772
rect 41244 9156 41300 9166
rect 41244 8818 41300 9100
rect 41244 8766 41246 8818
rect 41298 8766 41300 8818
rect 41244 8754 41300 8766
rect 41468 9044 41524 9054
rect 41468 8930 41524 8988
rect 41692 9042 41748 10108
rect 41916 10052 41972 10062
rect 41916 9826 41972 9996
rect 41916 9774 41918 9826
rect 41970 9774 41972 9826
rect 41916 9762 41972 9774
rect 42700 9940 42756 9950
rect 42812 9940 42868 10444
rect 43260 10434 43316 10444
rect 42756 9884 42868 9940
rect 42700 9604 42756 9884
rect 42700 9266 42756 9548
rect 43372 9380 43428 10668
rect 43820 10052 43876 20412
rect 44156 20244 44212 20254
rect 44156 20018 44212 20188
rect 44716 20130 44772 20524
rect 44828 20514 44884 20524
rect 45052 20468 45108 21084
rect 44716 20078 44718 20130
rect 44770 20078 44772 20130
rect 44716 20066 44772 20078
rect 44940 20412 45108 20468
rect 44156 19966 44158 20018
rect 44210 19966 44212 20018
rect 44156 19954 44212 19966
rect 44828 16212 44884 16222
rect 44828 16118 44884 16156
rect 44492 15988 44548 15998
rect 43932 15876 43988 15886
rect 43932 12964 43988 15820
rect 44044 15764 44100 15774
rect 44044 15314 44100 15708
rect 44492 15538 44548 15932
rect 44492 15486 44494 15538
rect 44546 15486 44548 15538
rect 44492 15474 44548 15486
rect 44604 15428 44660 15438
rect 44604 15334 44660 15372
rect 44044 15262 44046 15314
rect 44098 15262 44100 15314
rect 44044 15250 44100 15262
rect 44380 15204 44436 15242
rect 44380 15138 44436 15148
rect 43932 12962 44548 12964
rect 43932 12910 43934 12962
rect 43986 12910 44548 12962
rect 43932 12908 44548 12910
rect 43932 12898 43988 12908
rect 44492 12066 44548 12908
rect 44492 12014 44494 12066
rect 44546 12014 44548 12066
rect 44492 12002 44548 12014
rect 44828 11732 44884 11742
rect 44156 10948 44212 10958
rect 43820 9996 43988 10052
rect 43596 9716 43652 9726
rect 43596 9622 43652 9660
rect 42700 9214 42702 9266
rect 42754 9214 42756 9266
rect 42700 9202 42756 9214
rect 43260 9324 43428 9380
rect 41692 8990 41694 9042
rect 41746 8990 41748 9042
rect 41692 8978 41748 8990
rect 41916 9156 41972 9166
rect 41468 8878 41470 8930
rect 41522 8878 41524 8930
rect 41468 8370 41524 8878
rect 41468 8318 41470 8370
rect 41522 8318 41524 8370
rect 41468 8306 41524 8318
rect 41020 8206 41022 8258
rect 41074 8206 41076 8258
rect 41020 8194 41076 8206
rect 41804 8146 41860 8158
rect 41804 8094 41806 8146
rect 41858 8094 41860 8146
rect 41804 7924 41860 8094
rect 41916 8146 41972 9100
rect 43036 9042 43092 9054
rect 43036 8990 43038 9042
rect 43090 8990 43092 9042
rect 42812 8932 42868 8942
rect 41916 8094 41918 8146
rect 41970 8094 41972 8146
rect 41916 8082 41972 8094
rect 42252 8596 42308 8606
rect 42140 8036 42196 8046
rect 41804 7858 41860 7868
rect 42028 8034 42196 8036
rect 42028 7982 42142 8034
rect 42194 7982 42196 8034
rect 42028 7980 42196 7982
rect 41020 7700 41076 7710
rect 40908 7698 41076 7700
rect 40908 7646 41022 7698
rect 41074 7646 41076 7698
rect 40908 7644 41076 7646
rect 40908 7252 40964 7644
rect 41020 7634 41076 7644
rect 42028 7364 42084 7980
rect 42140 7970 42196 7980
rect 42140 7588 42196 7598
rect 42252 7588 42308 8540
rect 42476 8034 42532 8046
rect 42476 7982 42478 8034
rect 42530 7982 42532 8034
rect 42476 7924 42532 7982
rect 42476 7858 42532 7868
rect 42364 7700 42420 7710
rect 42364 7698 42756 7700
rect 42364 7646 42366 7698
rect 42418 7646 42756 7698
rect 42364 7644 42756 7646
rect 42364 7634 42420 7644
rect 42140 7586 42308 7588
rect 42140 7534 42142 7586
rect 42194 7534 42308 7586
rect 42140 7532 42308 7534
rect 42140 7522 42196 7532
rect 42588 7474 42644 7486
rect 42588 7422 42590 7474
rect 42642 7422 42644 7474
rect 42028 7308 42196 7364
rect 40348 7196 40964 7252
rect 40572 5234 40628 7196
rect 42140 6916 42196 7308
rect 42252 7252 42308 7262
rect 42252 7250 42420 7252
rect 42252 7198 42254 7250
rect 42306 7198 42420 7250
rect 42252 7196 42420 7198
rect 42252 7186 42308 7196
rect 42252 6916 42308 6926
rect 42140 6914 42308 6916
rect 42140 6862 42254 6914
rect 42306 6862 42308 6914
rect 42140 6860 42308 6862
rect 42028 6804 42084 6814
rect 42028 6802 42196 6804
rect 42028 6750 42030 6802
rect 42082 6750 42196 6802
rect 42028 6748 42196 6750
rect 42028 6738 42084 6748
rect 41804 6580 41860 6590
rect 41804 6486 41860 6524
rect 42028 6580 42084 6590
rect 40572 5182 40574 5234
rect 40626 5182 40628 5234
rect 39788 5068 40180 5124
rect 38892 5010 38948 5022
rect 38892 4958 38894 5010
rect 38946 4958 38948 5010
rect 37436 4900 37492 4910
rect 37436 4898 37716 4900
rect 37436 4846 37438 4898
rect 37490 4846 37716 4898
rect 37436 4844 37716 4846
rect 37436 4834 37492 4844
rect 37100 4610 37156 4620
rect 33180 4386 33236 4396
rect 33852 4452 33908 4462
rect 33852 4358 33908 4396
rect 33068 4340 33124 4350
rect 32956 4338 33124 4340
rect 32956 4286 33070 4338
rect 33122 4286 33124 4338
rect 32956 4284 33124 4286
rect 33068 4274 33124 4284
rect 36988 4338 37044 4508
rect 37660 4450 37716 4844
rect 37660 4398 37662 4450
rect 37714 4398 37716 4450
rect 37660 4386 37716 4398
rect 36988 4286 36990 4338
rect 37042 4286 37044 4338
rect 36988 4274 37044 4286
rect 32172 4174 32174 4226
rect 32226 4174 32228 4226
rect 32172 4162 32228 4174
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 38892 3780 38948 4958
rect 38892 3714 38948 3724
rect 39788 4898 39844 4910
rect 39788 4846 39790 4898
rect 39842 4846 39844 4898
rect 39788 4226 39844 4846
rect 39788 4174 39790 4226
rect 39842 4174 39844 4226
rect 39788 3780 39844 4174
rect 39788 3714 39844 3724
rect 29820 3668 29876 3678
rect 29036 3666 29316 3668
rect 29036 3614 29038 3666
rect 29090 3614 29316 3666
rect 29036 3612 29316 3614
rect 29596 3666 29876 3668
rect 29596 3614 29822 3666
rect 29874 3614 29876 3666
rect 29596 3612 29876 3614
rect 29036 3602 29092 3612
rect 11900 3502 11902 3554
rect 11954 3502 11956 3554
rect 11900 3490 11956 3502
rect 16156 3332 16212 3342
rect 16156 800 16212 3276
rect 16940 3332 16996 3342
rect 20860 3332 20916 3342
rect 25340 3332 25396 3342
rect 16940 3238 16996 3276
rect 20636 3330 20916 3332
rect 20636 3278 20862 3330
rect 20914 3278 20916 3330
rect 20636 3276 20916 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20636 800 20692 3276
rect 20860 3266 20916 3276
rect 25116 3330 25396 3332
rect 25116 3278 25342 3330
rect 25394 3278 25396 3330
rect 25116 3276 25396 3278
rect 25116 800 25172 3276
rect 25340 3266 25396 3276
rect 29596 800 29652 3612
rect 29820 3602 29876 3612
rect 34076 3668 34132 3678
rect 34076 800 34132 3612
rect 36988 3668 37044 3678
rect 40124 3668 40180 5068
rect 40236 4564 40292 4574
rect 40236 4470 40292 4508
rect 40572 4564 40628 5182
rect 41692 6132 41748 6142
rect 40572 4498 40628 4508
rect 41020 4564 41076 4574
rect 41020 4338 41076 4508
rect 41692 4450 41748 6076
rect 42028 6018 42084 6524
rect 42028 5966 42030 6018
rect 42082 5966 42084 6018
rect 42028 5954 42084 5966
rect 41804 5684 41860 5694
rect 42140 5684 42196 6748
rect 42252 5908 42308 6860
rect 42364 6132 42420 7196
rect 42364 6066 42420 6076
rect 42476 6692 42532 6702
rect 42364 5908 42420 5918
rect 42252 5906 42420 5908
rect 42252 5854 42366 5906
rect 42418 5854 42420 5906
rect 42252 5852 42420 5854
rect 42476 5908 42532 6636
rect 42588 6132 42644 7422
rect 42700 6916 42756 7644
rect 42812 7586 42868 8876
rect 43036 8484 43092 8990
rect 43036 8418 43092 8428
rect 42812 7534 42814 7586
rect 42866 7534 42868 7586
rect 42812 7522 42868 7534
rect 42924 6916 42980 6926
rect 42700 6914 42980 6916
rect 42700 6862 42926 6914
rect 42978 6862 42980 6914
rect 42700 6860 42980 6862
rect 42924 6850 42980 6860
rect 42700 6132 42756 6142
rect 42588 6130 42756 6132
rect 42588 6078 42702 6130
rect 42754 6078 42756 6130
rect 42588 6076 42756 6078
rect 42700 6066 42756 6076
rect 42588 5908 42644 5918
rect 42476 5906 42644 5908
rect 42476 5854 42590 5906
rect 42642 5854 42644 5906
rect 42476 5852 42644 5854
rect 42364 5842 42420 5852
rect 42588 5842 42644 5852
rect 43260 5908 43316 9324
rect 43372 9156 43428 9166
rect 43372 8596 43428 9100
rect 43372 7698 43428 8540
rect 43372 7646 43374 7698
rect 43426 7646 43428 7698
rect 43372 7634 43428 7646
rect 43260 5842 43316 5852
rect 41804 5682 42196 5684
rect 41804 5630 41806 5682
rect 41858 5630 42196 5682
rect 41804 5628 42196 5630
rect 41804 5618 41860 5628
rect 42140 5124 42196 5628
rect 42140 5058 42196 5068
rect 43820 5124 43876 5134
rect 41692 4398 41694 4450
rect 41746 4398 41748 4450
rect 41692 4386 41748 4398
rect 41020 4286 41022 4338
rect 41074 4286 41076 4338
rect 41020 4274 41076 4286
rect 43820 4226 43876 5068
rect 43932 5012 43988 9996
rect 44044 7700 44100 7710
rect 44044 7364 44100 7644
rect 44044 7298 44100 7308
rect 44044 5012 44100 5022
rect 43932 4956 44044 5012
rect 44044 4946 44100 4956
rect 43820 4174 43822 4226
rect 43874 4174 43876 4226
rect 43820 4162 43876 4174
rect 40236 3668 40292 3678
rect 40124 3666 40292 3668
rect 40124 3614 40238 3666
rect 40290 3614 40292 3666
rect 40124 3612 40292 3614
rect 36988 3574 37044 3612
rect 40236 3602 40292 3612
rect 35532 3556 35588 3566
rect 35532 3462 35588 3500
rect 35980 3556 36036 3566
rect 35980 3462 36036 3500
rect 38556 3444 38612 3454
rect 38556 800 38612 3388
rect 39340 3444 39396 3482
rect 39340 3378 39396 3388
rect 39788 3444 39844 3482
rect 43148 3444 43204 3454
rect 43596 3444 43652 3454
rect 39788 3378 39844 3388
rect 43036 3442 43652 3444
rect 43036 3390 43150 3442
rect 43202 3390 43598 3442
rect 43650 3390 43652 3442
rect 43036 3388 43652 3390
rect 43036 800 43092 3388
rect 43148 3378 43204 3388
rect 43596 3378 43652 3388
rect 43932 3444 43988 3454
rect 44156 3444 44212 10892
rect 44268 10610 44324 10622
rect 44268 10558 44270 10610
rect 44322 10558 44324 10610
rect 44268 9828 44324 10558
rect 44492 10610 44548 10622
rect 44492 10558 44494 10610
rect 44546 10558 44548 10610
rect 44268 9762 44324 9772
rect 44380 10498 44436 10510
rect 44380 10446 44382 10498
rect 44434 10446 44436 10498
rect 44268 9604 44324 9614
rect 44268 9510 44324 9548
rect 44380 8932 44436 10446
rect 44492 10164 44548 10558
rect 44828 10610 44884 11676
rect 44828 10558 44830 10610
rect 44882 10558 44884 10610
rect 44828 10546 44884 10558
rect 44492 10098 44548 10108
rect 44380 8866 44436 8876
rect 44828 8372 44884 8382
rect 44268 7700 44324 7710
rect 44268 7698 44772 7700
rect 44268 7646 44270 7698
rect 44322 7646 44772 7698
rect 44268 7644 44772 7646
rect 44268 7634 44324 7644
rect 44716 5236 44772 7644
rect 44828 7474 44884 8316
rect 44828 7422 44830 7474
rect 44882 7422 44884 7474
rect 44828 7410 44884 7422
rect 44940 6132 44996 20412
rect 45052 18340 45108 18350
rect 45052 18246 45108 18284
rect 45164 15148 45220 21308
rect 45276 20692 45332 21420
rect 45388 21410 45444 21420
rect 45388 20916 45444 20926
rect 45500 20916 45556 21868
rect 46396 21812 46452 21822
rect 46396 21718 46452 21756
rect 45836 21588 45892 21598
rect 45836 21494 45892 21532
rect 45388 20914 45556 20916
rect 45388 20862 45390 20914
rect 45442 20862 45556 20914
rect 45388 20860 45556 20862
rect 45724 21028 45780 21038
rect 45388 20850 45444 20860
rect 45276 20636 45444 20692
rect 45052 15092 45220 15148
rect 45388 15148 45444 20636
rect 45500 20244 45556 20254
rect 45500 19906 45556 20188
rect 45500 19854 45502 19906
rect 45554 19854 45556 19906
rect 45500 19842 45556 19854
rect 45612 19236 45668 19246
rect 45500 18564 45556 18574
rect 45500 18470 45556 18508
rect 45388 15092 45556 15148
rect 45052 10948 45108 15092
rect 45388 12516 45444 12526
rect 45388 12402 45444 12460
rect 45388 12350 45390 12402
rect 45442 12350 45444 12402
rect 45388 12338 45444 12350
rect 45500 11788 45556 15092
rect 45388 11732 45556 11788
rect 45612 12740 45668 19180
rect 45724 14420 45780 20972
rect 46508 21028 46564 28700
rect 46956 28642 47012 29260
rect 47068 29250 47124 29260
rect 46956 28590 46958 28642
rect 47010 28590 47012 28642
rect 46956 28578 47012 28590
rect 47068 28756 47124 28766
rect 47068 28642 47124 28700
rect 47068 28590 47070 28642
rect 47122 28590 47124 28642
rect 47068 28578 47124 28590
rect 47180 28532 47236 28542
rect 47180 28438 47236 28476
rect 47404 28084 47460 34636
rect 48188 34692 48244 34702
rect 48188 34018 48244 34636
rect 48188 33966 48190 34018
rect 48242 33966 48244 34018
rect 48188 33954 48244 33966
rect 47740 31890 47796 31902
rect 47740 31838 47742 31890
rect 47794 31838 47796 31890
rect 47740 30324 47796 31838
rect 47964 31556 48020 31566
rect 47964 30994 48020 31500
rect 48188 31332 48244 31342
rect 48188 31218 48244 31276
rect 48188 31166 48190 31218
rect 48242 31166 48244 31218
rect 48188 31154 48244 31166
rect 47964 30942 47966 30994
rect 48018 30942 48020 30994
rect 47964 30930 48020 30942
rect 47740 28532 47796 30268
rect 48300 28868 48356 40908
rect 48412 40898 48468 40908
rect 48636 37268 48692 37278
rect 48748 37268 48804 42700
rect 49308 42420 49364 42430
rect 48860 41972 48916 41982
rect 48860 41878 48916 41916
rect 49308 41970 49364 42364
rect 49308 41918 49310 41970
rect 49362 41918 49364 41970
rect 49308 41906 49364 41918
rect 49644 41748 49700 41758
rect 49084 41746 49700 41748
rect 49084 41694 49646 41746
rect 49698 41694 49700 41746
rect 49084 41692 49700 41694
rect 49084 41298 49140 41692
rect 49644 41682 49700 41692
rect 49084 41246 49086 41298
rect 49138 41246 49140 41298
rect 49084 41234 49140 41246
rect 49196 41188 49252 41198
rect 49196 41094 49252 41132
rect 49756 41188 49812 44380
rect 49980 44098 50036 44110
rect 49980 44046 49982 44098
rect 50034 44046 50036 44098
rect 49980 43764 50036 44046
rect 49980 42530 50036 43708
rect 49980 42478 49982 42530
rect 50034 42478 50036 42530
rect 49868 42420 49924 42430
rect 49868 42194 49924 42364
rect 49868 42142 49870 42194
rect 49922 42142 49924 42194
rect 49868 42130 49924 42142
rect 49980 41972 50036 42478
rect 50204 42420 50260 45836
rect 50316 43764 50372 46508
rect 50556 45500 50820 45510
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50556 45434 50820 45444
rect 51212 45332 51268 47068
rect 50988 45276 51268 45332
rect 50988 44324 51044 45276
rect 51100 45106 51156 45118
rect 51100 45054 51102 45106
rect 51154 45054 51156 45106
rect 51100 44436 51156 45054
rect 51100 44380 51380 44436
rect 50988 44268 51268 44324
rect 50540 44212 50596 44222
rect 50540 44118 50596 44156
rect 50876 44098 50932 44110
rect 50876 44046 50878 44098
rect 50930 44046 50932 44098
rect 50556 43932 50820 43942
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50556 43866 50820 43876
rect 50316 43538 50372 43708
rect 50876 43708 50932 44046
rect 50876 43652 51156 43708
rect 51100 43650 51156 43652
rect 51100 43598 51102 43650
rect 51154 43598 51156 43650
rect 51100 43586 51156 43598
rect 50316 43486 50318 43538
rect 50370 43486 50372 43538
rect 50316 43474 50372 43486
rect 50316 42420 50372 42430
rect 50204 42364 50316 42420
rect 49980 41906 50036 41916
rect 49868 41860 49924 41870
rect 49868 41766 49924 41804
rect 49756 41122 49812 41132
rect 49980 41186 50036 41198
rect 49980 41134 49982 41186
rect 50034 41134 50036 41186
rect 48972 40962 49028 40974
rect 48972 40910 48974 40962
rect 49026 40910 49028 40962
rect 48860 39506 48916 39518
rect 48860 39454 48862 39506
rect 48914 39454 48916 39506
rect 48860 39172 48916 39454
rect 48860 39106 48916 39116
rect 48972 37380 49028 40910
rect 49644 39620 49700 39630
rect 49532 39396 49588 39406
rect 49308 39284 49364 39294
rect 49308 37490 49364 39228
rect 49308 37438 49310 37490
rect 49362 37438 49364 37490
rect 49084 37380 49140 37390
rect 48636 37266 48804 37268
rect 48636 37214 48638 37266
rect 48690 37214 48804 37266
rect 48636 37212 48804 37214
rect 48860 37378 49140 37380
rect 48860 37326 49086 37378
rect 49138 37326 49140 37378
rect 48860 37324 49140 37326
rect 48636 37044 48692 37212
rect 48636 36978 48692 36988
rect 48860 34468 48916 37324
rect 49084 37314 49140 37324
rect 49196 37156 49252 37166
rect 49196 37062 49252 37100
rect 49308 36932 49364 37438
rect 48972 36876 49364 36932
rect 48972 36594 49028 36876
rect 48972 36542 48974 36594
rect 49026 36542 49028 36594
rect 48972 36530 49028 36542
rect 49420 35698 49476 35710
rect 49420 35646 49422 35698
rect 49474 35646 49476 35698
rect 49084 35588 49140 35598
rect 49420 35588 49476 35646
rect 49140 35532 49476 35588
rect 49084 35494 49140 35532
rect 49308 34692 49364 34702
rect 48860 34412 49140 34468
rect 49084 34354 49140 34412
rect 49084 34302 49086 34354
rect 49138 34302 49140 34354
rect 48748 34130 48804 34142
rect 48748 34078 48750 34130
rect 48802 34078 48804 34130
rect 48748 33572 48804 34078
rect 48412 33516 48804 33572
rect 48412 33460 48468 33516
rect 49084 33460 49140 34302
rect 49308 34354 49364 34636
rect 49308 34302 49310 34354
rect 49362 34302 49364 34354
rect 49308 34290 49364 34302
rect 49308 34132 49364 34142
rect 49196 34018 49252 34030
rect 49196 33966 49198 34018
rect 49250 33966 49252 34018
rect 49196 33684 49252 33966
rect 49196 33618 49252 33628
rect 49084 33404 49252 33460
rect 48412 33366 48468 33404
rect 49084 31668 49140 31678
rect 49084 31574 49140 31612
rect 48748 31556 48804 31566
rect 48748 31462 48804 31500
rect 49196 31332 49252 33404
rect 49308 31780 49364 34076
rect 49308 31714 49364 31724
rect 49420 31892 49476 31902
rect 49196 31218 49252 31276
rect 49196 31166 49198 31218
rect 49250 31166 49252 31218
rect 49196 31154 49252 31166
rect 49420 31218 49476 31836
rect 49420 31166 49422 31218
rect 49474 31166 49476 31218
rect 49420 31154 49476 31166
rect 48748 30996 48804 31006
rect 48748 30902 48804 30940
rect 48972 30882 49028 30894
rect 48972 30830 48974 30882
rect 49026 30830 49028 30882
rect 48972 30772 49028 30830
rect 48972 30706 49028 30716
rect 49308 30882 49364 30894
rect 49308 30830 49310 30882
rect 49362 30830 49364 30882
rect 49308 30436 49364 30830
rect 49308 30370 49364 30380
rect 48300 28802 48356 28812
rect 48076 28644 48132 28654
rect 48076 28550 48132 28588
rect 47740 28466 47796 28476
rect 48748 28530 48804 28542
rect 48748 28478 48750 28530
rect 48802 28478 48804 28530
rect 47404 28018 47460 28028
rect 47628 28418 47684 28430
rect 47628 28366 47630 28418
rect 47682 28366 47684 28418
rect 47628 26908 47684 28366
rect 48300 28084 48356 28094
rect 48748 28084 48804 28478
rect 49532 28308 49588 39340
rect 49644 38836 49700 39564
rect 49644 38770 49700 38780
rect 49980 38668 50036 41134
rect 50316 40404 50372 42364
rect 50556 42364 50820 42374
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50556 42298 50820 42308
rect 50428 41972 50484 41982
rect 50428 41878 50484 41916
rect 51100 41860 51156 41870
rect 51100 41766 51156 41804
rect 50556 40796 50820 40806
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50556 40730 50820 40740
rect 51212 40628 51268 44268
rect 51324 43708 51380 44380
rect 51548 43708 51604 47630
rect 51660 47234 51716 47246
rect 51660 47182 51662 47234
rect 51714 47182 51716 47234
rect 51660 46676 51716 47182
rect 51660 46610 51716 46620
rect 53004 46228 53060 47966
rect 53228 46900 53284 46910
rect 53228 46562 53284 46844
rect 53228 46510 53230 46562
rect 53282 46510 53284 46562
rect 53228 46498 53284 46510
rect 53004 46162 53060 46172
rect 53004 44882 53060 44894
rect 53004 44830 53006 44882
rect 53058 44830 53060 44882
rect 51324 43652 51492 43708
rect 51548 43652 51828 43708
rect 50764 40572 51268 40628
rect 50316 40348 50484 40404
rect 50316 39618 50372 39630
rect 50316 39566 50318 39618
rect 50370 39566 50372 39618
rect 50204 39396 50260 39406
rect 50316 39396 50372 39566
rect 50428 39508 50484 40348
rect 50428 39442 50484 39452
rect 50652 40402 50708 40414
rect 50652 40350 50654 40402
rect 50706 40350 50708 40402
rect 50260 39340 50372 39396
rect 50652 39396 50708 40350
rect 50764 39620 50820 40572
rect 50764 39526 50820 39564
rect 50876 39620 50932 39630
rect 51324 39620 51380 39630
rect 50876 39618 51380 39620
rect 50876 39566 50878 39618
rect 50930 39566 51326 39618
rect 51378 39566 51380 39618
rect 50876 39564 51380 39566
rect 51436 39620 51492 43652
rect 51772 39732 51828 43652
rect 53004 43540 53060 44830
rect 53004 43474 53060 43484
rect 53228 43428 53284 43438
rect 53228 43334 53284 43372
rect 53228 41858 53284 41870
rect 53228 41806 53230 41858
rect 53282 41806 53284 41858
rect 51884 41298 51940 41310
rect 51884 41246 51886 41298
rect 51938 41246 51940 41298
rect 51884 40852 51940 41246
rect 53228 41188 53284 41806
rect 53228 41122 53284 41132
rect 51884 40786 51940 40796
rect 53004 40178 53060 40190
rect 53004 40126 53006 40178
rect 53058 40126 53060 40178
rect 51772 39676 51940 39732
rect 51436 39564 51828 39620
rect 50876 39554 50932 39564
rect 51324 39554 51380 39564
rect 50988 39396 51044 39406
rect 50204 39302 50260 39340
rect 50652 39330 50708 39340
rect 50876 39394 51044 39396
rect 50876 39342 50990 39394
rect 51042 39342 51044 39394
rect 50876 39340 51044 39342
rect 50556 39228 50820 39238
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50556 39162 50820 39172
rect 49644 38612 50036 38668
rect 50428 38836 50484 38846
rect 49644 31556 49700 38612
rect 50428 37266 50484 38780
rect 50556 37660 50820 37670
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50556 37594 50820 37604
rect 50428 37214 50430 37266
rect 50482 37214 50484 37266
rect 50092 36482 50148 36494
rect 50092 36430 50094 36482
rect 50146 36430 50148 36482
rect 49756 35812 49812 35822
rect 49756 34242 49812 35756
rect 49756 34190 49758 34242
rect 49810 34190 49812 34242
rect 49756 33572 49812 34190
rect 49980 34132 50036 34142
rect 50092 34132 50148 36430
rect 50036 34076 50148 34132
rect 50316 34132 50372 34142
rect 50428 34132 50484 37214
rect 50876 36820 50932 39340
rect 50988 39330 51044 39340
rect 51436 39394 51492 39406
rect 51436 39342 51438 39394
rect 51490 39342 51492 39394
rect 51436 39060 51492 39342
rect 51548 39396 51604 39406
rect 51548 39302 51604 39340
rect 51100 39004 51492 39060
rect 51100 38946 51156 39004
rect 51100 38894 51102 38946
rect 51154 38894 51156 38946
rect 51100 38882 51156 38894
rect 51100 37156 51156 37166
rect 51100 37154 51268 37156
rect 51100 37102 51102 37154
rect 51154 37102 51268 37154
rect 51100 37100 51268 37102
rect 51100 37090 51156 37100
rect 50540 36764 50932 36820
rect 50988 37044 51044 37054
rect 50540 36482 50596 36764
rect 50988 36708 51044 36988
rect 50876 36652 51044 36708
rect 50540 36430 50542 36482
rect 50594 36430 50596 36482
rect 50540 36260 50596 36430
rect 50764 36484 50820 36494
rect 50876 36484 50932 36652
rect 51212 36594 51268 37100
rect 51212 36542 51214 36594
rect 51266 36542 51268 36594
rect 51212 36530 51268 36542
rect 50764 36482 50932 36484
rect 50764 36430 50766 36482
rect 50818 36430 50932 36482
rect 50764 36428 50932 36430
rect 50764 36418 50820 36428
rect 50652 36372 50708 36382
rect 50652 36278 50708 36316
rect 51100 36372 51156 36382
rect 51100 36278 51156 36316
rect 50540 36194 50596 36204
rect 50876 36260 50932 36270
rect 50556 36092 50820 36102
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50556 36026 50820 36036
rect 50652 35698 50708 35710
rect 50652 35646 50654 35698
rect 50706 35646 50708 35698
rect 50652 34692 50708 35646
rect 50652 34626 50708 34636
rect 50556 34524 50820 34534
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50556 34458 50820 34468
rect 50316 34130 50484 34132
rect 50316 34078 50318 34130
rect 50370 34078 50484 34130
rect 50316 34076 50484 34078
rect 49980 34066 50036 34076
rect 50316 34066 50372 34076
rect 49868 34020 49924 34030
rect 49868 33926 49924 33964
rect 49980 33906 50036 33918
rect 49980 33854 49982 33906
rect 50034 33854 50036 33906
rect 49980 33572 50036 33854
rect 50540 33908 50596 33918
rect 49980 33516 50260 33572
rect 49756 33506 49812 33516
rect 50204 33460 50260 33516
rect 50428 33460 50484 33470
rect 50204 33458 50484 33460
rect 50204 33406 50430 33458
rect 50482 33406 50484 33458
rect 50204 33404 50484 33406
rect 50428 33394 50484 33404
rect 49868 33346 49924 33358
rect 49868 33294 49870 33346
rect 49922 33294 49924 33346
rect 49868 32788 49924 33294
rect 50540 33346 50596 33852
rect 50540 33294 50542 33346
rect 50594 33294 50596 33346
rect 50540 33282 50596 33294
rect 50316 33124 50372 33134
rect 50876 33124 50932 36204
rect 51324 36258 51380 36270
rect 51324 36206 51326 36258
rect 51378 36206 51380 36258
rect 51324 35812 51380 36206
rect 51324 35746 51380 35756
rect 51100 34020 51156 34030
rect 51100 33926 51156 33964
rect 51772 34020 51828 39564
rect 51884 37044 51940 39676
rect 52108 39508 52164 39518
rect 52108 39414 52164 39452
rect 53004 38164 53060 40126
rect 53228 39620 53284 39630
rect 53228 38722 53284 39564
rect 53228 38670 53230 38722
rect 53282 38670 53284 38722
rect 53228 38658 53284 38670
rect 53004 38098 53060 38108
rect 51884 36978 51940 36988
rect 53228 37154 53284 37166
rect 53228 37102 53230 37154
rect 53282 37102 53284 37154
rect 53228 37044 53284 37102
rect 53228 36978 53284 36988
rect 53004 35476 53060 35486
rect 53004 35382 53060 35420
rect 51772 33954 51828 33964
rect 53228 34020 53284 34030
rect 53228 33926 53284 33964
rect 50316 33122 50932 33124
rect 50316 33070 50318 33122
rect 50370 33070 50932 33122
rect 50316 33068 50932 33070
rect 51212 33572 51268 33582
rect 50316 33058 50372 33068
rect 49868 32722 49924 32732
rect 49980 31778 50036 31790
rect 49980 31726 49982 31778
rect 50034 31726 50036 31778
rect 49756 31556 49812 31566
rect 49644 31500 49756 31556
rect 49756 31490 49812 31500
rect 49980 31220 50036 31726
rect 50428 31780 50484 33068
rect 50556 32956 50820 32966
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50556 32890 50820 32900
rect 51100 32562 51156 32574
rect 51100 32510 51102 32562
rect 51154 32510 51156 32562
rect 50428 31686 50484 31724
rect 50540 31780 50596 31790
rect 50988 31780 51044 31790
rect 50540 31778 51044 31780
rect 50540 31726 50542 31778
rect 50594 31726 50990 31778
rect 51042 31726 51044 31778
rect 50540 31724 51044 31726
rect 50540 31714 50596 31724
rect 50988 31714 51044 31724
rect 51100 31780 51156 32510
rect 51100 31714 51156 31724
rect 51212 31666 51268 33516
rect 53004 32788 53060 32798
rect 53004 32450 53060 32732
rect 53004 32398 53006 32450
rect 53058 32398 53060 32450
rect 53004 32386 53060 32398
rect 51212 31614 51214 31666
rect 51266 31614 51268 31666
rect 50652 31556 50708 31594
rect 50652 31490 50708 31500
rect 51100 31554 51156 31566
rect 51100 31502 51102 31554
rect 51154 31502 51156 31554
rect 50556 31388 50820 31398
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50556 31322 50820 31332
rect 49980 31154 50036 31164
rect 51100 31106 51156 31502
rect 51100 31054 51102 31106
rect 51154 31054 51156 31106
rect 51100 31042 51156 31054
rect 50428 30994 50484 31006
rect 50428 30942 50430 30994
rect 50482 30942 50484 30994
rect 50428 30548 50484 30942
rect 50316 30492 50484 30548
rect 50204 30436 50260 30446
rect 50204 30342 50260 30380
rect 50316 30100 50372 30492
rect 51212 30436 51268 31614
rect 50652 30380 51268 30436
rect 53116 31780 53172 31790
rect 50428 30324 50484 30334
rect 50428 30230 50484 30268
rect 50540 30210 50596 30222
rect 50540 30158 50542 30210
rect 50594 30158 50596 30210
rect 50540 30100 50596 30158
rect 50652 30100 50708 30380
rect 50316 30044 50484 30100
rect 50540 30044 50708 30100
rect 51100 30212 51156 30222
rect 49532 28242 49588 28252
rect 50428 29426 50484 30044
rect 50556 29820 50820 29830
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50556 29754 50820 29764
rect 51100 29538 51156 30156
rect 52220 30100 52276 30110
rect 52220 30006 52276 30044
rect 52892 29988 52948 29998
rect 51100 29486 51102 29538
rect 51154 29486 51156 29538
rect 51100 29474 51156 29486
rect 52332 29986 52948 29988
rect 52332 29934 52894 29986
rect 52946 29934 52948 29986
rect 52332 29932 52948 29934
rect 50428 29374 50430 29426
rect 50482 29374 50484 29426
rect 50428 28644 50484 29374
rect 48860 28084 48916 28094
rect 48748 28082 48916 28084
rect 48748 28030 48862 28082
rect 48914 28030 48916 28082
rect 48748 28028 48916 28030
rect 48300 27990 48356 28028
rect 48860 28018 48916 28028
rect 48972 28084 49028 28094
rect 48972 27990 49028 28028
rect 48748 27634 48804 27646
rect 48748 27582 48750 27634
rect 48802 27582 48804 27634
rect 48748 26908 48804 27582
rect 47516 26852 47684 26908
rect 48076 26852 48804 26908
rect 49644 26964 49700 26974
rect 47068 24052 47124 24062
rect 47068 23958 47124 23996
rect 46732 23714 46788 23726
rect 46732 23662 46734 23714
rect 46786 23662 46788 23714
rect 46732 23604 46788 23662
rect 46732 23538 46788 23548
rect 46508 20962 46564 20972
rect 46620 23492 46676 23502
rect 46620 22036 46676 23436
rect 45948 20804 46004 20814
rect 45948 20710 46004 20748
rect 46508 20804 46564 20814
rect 46508 20710 46564 20748
rect 45836 20580 45892 20590
rect 46620 20580 46676 21980
rect 47292 21588 47348 21598
rect 47292 21494 47348 21532
rect 45836 19012 45892 20524
rect 46508 20524 46676 20580
rect 46732 21474 46788 21486
rect 46732 21422 46734 21474
rect 46786 21422 46788 21474
rect 46396 20244 46452 20254
rect 46284 20020 46340 20030
rect 46172 20018 46340 20020
rect 46172 19966 46286 20018
rect 46338 19966 46340 20018
rect 46172 19964 46340 19966
rect 45948 19908 46004 19918
rect 45948 19346 46004 19852
rect 45948 19294 45950 19346
rect 46002 19294 46004 19346
rect 45948 19236 46004 19294
rect 45948 19170 46004 19180
rect 46060 19796 46116 19806
rect 45836 18956 46004 19012
rect 45836 18562 45892 18574
rect 45836 18510 45838 18562
rect 45890 18510 45892 18562
rect 45836 18452 45892 18510
rect 45836 18386 45892 18396
rect 45724 14354 45780 14364
rect 45836 15540 45892 15550
rect 45388 11284 45444 11732
rect 45388 11218 45444 11228
rect 45612 11284 45668 12684
rect 45724 12516 45780 12526
rect 45836 12516 45892 15484
rect 45948 12964 46004 18956
rect 46060 14980 46116 19740
rect 46172 18564 46228 19964
rect 46284 19954 46340 19964
rect 46284 19236 46340 19246
rect 46284 19142 46340 19180
rect 46172 18498 46228 18508
rect 46172 18340 46228 18350
rect 46172 18246 46228 18284
rect 46396 15540 46452 20188
rect 46508 18228 46564 20524
rect 46620 19236 46676 19246
rect 46620 19122 46676 19180
rect 46620 19070 46622 19122
rect 46674 19070 46676 19122
rect 46620 19058 46676 19070
rect 46732 19012 46788 21422
rect 46956 20580 47012 20590
rect 46956 20486 47012 20524
rect 47404 20578 47460 20590
rect 47404 20526 47406 20578
rect 47458 20526 47460 20578
rect 47404 20244 47460 20526
rect 47404 20178 47460 20188
rect 46844 19906 46900 19918
rect 46844 19854 46846 19906
rect 46898 19854 46900 19906
rect 46844 19796 46900 19854
rect 46844 19730 46900 19740
rect 46732 18946 46788 18956
rect 46732 18450 46788 18462
rect 46732 18398 46734 18450
rect 46786 18398 46788 18450
rect 46732 18340 46788 18398
rect 47180 18340 47236 18350
rect 46732 18338 47236 18340
rect 46732 18286 47182 18338
rect 47234 18286 47236 18338
rect 46732 18284 47236 18286
rect 46508 18172 46900 18228
rect 46732 15540 46788 15550
rect 46452 15538 46788 15540
rect 46452 15486 46734 15538
rect 46786 15486 46788 15538
rect 46452 15484 46788 15486
rect 46396 15446 46452 15484
rect 46732 15474 46788 15484
rect 46844 15148 46900 18172
rect 47180 17444 47236 18284
rect 47180 17378 47236 17388
rect 46956 15988 47012 15998
rect 46956 15894 47012 15932
rect 47068 15428 47124 15438
rect 47068 15204 47124 15372
rect 46060 14914 46116 14924
rect 46396 15092 46452 15102
rect 46844 15092 47012 15148
rect 47068 15138 47124 15148
rect 47516 15148 47572 26852
rect 47964 26178 48020 26190
rect 47964 26126 47966 26178
rect 48018 26126 48020 26178
rect 47740 25508 47796 25518
rect 47740 25414 47796 25452
rect 47964 25396 48020 26126
rect 47964 25330 48020 25340
rect 48076 25282 48132 26852
rect 49420 26290 49476 26302
rect 49420 26238 49422 26290
rect 49474 26238 49476 26290
rect 49420 25508 49476 26238
rect 49644 26290 49700 26908
rect 49644 26238 49646 26290
rect 49698 26238 49700 26290
rect 49532 26180 49588 26190
rect 49532 26086 49588 26124
rect 49644 25956 49700 26238
rect 49420 25442 49476 25452
rect 49532 25900 49700 25956
rect 49868 26290 49924 26302
rect 49868 26238 49870 26290
rect 49922 26238 49924 26290
rect 48188 25396 48244 25406
rect 48188 25302 48244 25340
rect 48412 25394 48468 25406
rect 48412 25342 48414 25394
rect 48466 25342 48468 25394
rect 48076 25230 48078 25282
rect 48130 25230 48132 25282
rect 48076 25218 48132 25230
rect 48412 25284 48468 25342
rect 48412 25218 48468 25228
rect 48748 25394 48804 25406
rect 48748 25342 48750 25394
rect 48802 25342 48804 25394
rect 47628 23716 47684 23726
rect 48748 23716 48804 25342
rect 49084 25396 49140 25406
rect 49308 25396 49364 25406
rect 49084 25394 49252 25396
rect 49084 25342 49086 25394
rect 49138 25342 49252 25394
rect 49084 25340 49252 25342
rect 49084 25330 49140 25340
rect 48860 25284 48916 25294
rect 48860 25190 48916 25228
rect 49196 24948 49252 25340
rect 49308 25302 49364 25340
rect 49308 24948 49364 24958
rect 49196 24946 49364 24948
rect 49196 24894 49310 24946
rect 49362 24894 49364 24946
rect 49196 24892 49364 24894
rect 49308 24882 49364 24892
rect 49532 24946 49588 25900
rect 49868 25732 49924 26238
rect 49756 25676 49924 25732
rect 50428 26290 50484 28588
rect 50876 28754 50932 28766
rect 50876 28702 50878 28754
rect 50930 28702 50932 28754
rect 50556 28252 50820 28262
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50556 28186 50820 28196
rect 50876 26964 50932 28702
rect 50876 26898 50932 26908
rect 50556 26684 50820 26694
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50556 26618 50820 26628
rect 50428 26238 50430 26290
rect 50482 26238 50484 26290
rect 49756 25618 49812 25676
rect 49756 25566 49758 25618
rect 49810 25566 49812 25618
rect 49756 25554 49812 25566
rect 50092 25620 50148 25630
rect 49868 25506 49924 25518
rect 49868 25454 49870 25506
rect 49922 25454 49924 25506
rect 49644 25396 49700 25406
rect 49644 25394 49812 25396
rect 49644 25342 49646 25394
rect 49698 25342 49812 25394
rect 49644 25340 49812 25342
rect 49644 25330 49700 25340
rect 49532 24894 49534 24946
rect 49586 24894 49588 24946
rect 49532 24882 49588 24894
rect 49644 24722 49700 24734
rect 49644 24670 49646 24722
rect 49698 24670 49700 24722
rect 49084 24612 49140 24622
rect 49084 24518 49140 24556
rect 49644 24612 49700 24670
rect 49644 24546 49700 24556
rect 49756 24164 49812 25340
rect 49868 24946 49924 25454
rect 49868 24894 49870 24946
rect 49922 24894 49924 24946
rect 49868 24882 49924 24894
rect 49084 24108 49812 24164
rect 50092 24834 50148 25564
rect 50204 25396 50260 25406
rect 50260 25340 50372 25396
rect 50204 25302 50260 25340
rect 50092 24782 50094 24834
rect 50146 24782 50148 24834
rect 48748 23660 49028 23716
rect 47628 23622 47684 23660
rect 48300 23604 48356 23614
rect 48188 23492 48356 23548
rect 47964 23044 48020 23054
rect 47964 22950 48020 22988
rect 48076 22482 48132 22494
rect 48076 22430 48078 22482
rect 48130 22430 48132 22482
rect 47852 22148 47908 22158
rect 47628 21586 47684 21598
rect 47628 21534 47630 21586
rect 47682 21534 47684 21586
rect 47628 20244 47684 21534
rect 47628 20178 47684 20188
rect 47852 19236 47908 22092
rect 47964 21700 48020 21710
rect 47964 21606 48020 21644
rect 48076 20916 48132 22430
rect 48076 20850 48132 20860
rect 48188 19460 48244 23492
rect 48860 23380 48916 23390
rect 48636 23378 48916 23380
rect 48636 23326 48862 23378
rect 48914 23326 48916 23378
rect 48636 23324 48916 23326
rect 48636 21588 48692 23324
rect 48860 23314 48916 23324
rect 48748 23154 48804 23166
rect 48748 23102 48750 23154
rect 48802 23102 48804 23154
rect 48748 22372 48804 23102
rect 48860 22596 48916 22606
rect 48972 22596 49028 23660
rect 49084 23378 49140 24108
rect 50092 24052 50148 24782
rect 50204 24722 50260 24734
rect 50204 24670 50206 24722
rect 50258 24670 50260 24722
rect 50204 24612 50260 24670
rect 50204 24546 50260 24556
rect 49756 23996 50148 24052
rect 49084 23326 49086 23378
rect 49138 23326 49140 23378
rect 49084 23314 49140 23326
rect 49420 23716 49476 23726
rect 49308 23154 49364 23166
rect 49308 23102 49310 23154
rect 49362 23102 49364 23154
rect 49308 22932 49364 23102
rect 49308 22866 49364 22876
rect 48860 22594 49028 22596
rect 48860 22542 48862 22594
rect 48914 22542 49028 22594
rect 48860 22540 49028 22542
rect 48860 22530 48916 22540
rect 48972 22372 49028 22382
rect 49308 22372 49364 22382
rect 48748 22370 49028 22372
rect 48748 22318 48974 22370
rect 49026 22318 49028 22370
rect 48748 22316 49028 22318
rect 48748 21700 48804 22316
rect 48972 22306 49028 22316
rect 49084 22370 49364 22372
rect 49084 22318 49310 22370
rect 49362 22318 49364 22370
rect 49084 22316 49364 22318
rect 48860 22148 48916 22158
rect 48860 22054 48916 22092
rect 49084 21810 49140 22316
rect 49308 22306 49364 22316
rect 49420 22260 49476 23660
rect 49756 23266 49812 23996
rect 49756 23214 49758 23266
rect 49810 23214 49812 23266
rect 49756 23202 49812 23214
rect 49868 23154 49924 23166
rect 49868 23102 49870 23154
rect 49922 23102 49924 23154
rect 49532 23044 49588 23054
rect 49532 22950 49588 22988
rect 49868 22596 49924 23102
rect 50316 22820 50372 25340
rect 50428 23268 50484 26238
rect 50988 26180 51044 26190
rect 50988 25730 51044 26124
rect 50988 25678 50990 25730
rect 51042 25678 51044 25730
rect 50988 25666 51044 25678
rect 51100 26178 51156 26190
rect 51100 26126 51102 26178
rect 51154 26126 51156 26178
rect 51100 25618 51156 26126
rect 51100 25566 51102 25618
rect 51154 25566 51156 25618
rect 51100 25554 51156 25566
rect 51212 25282 51268 25294
rect 51212 25230 51214 25282
rect 51266 25230 51268 25282
rect 50556 25116 50820 25126
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50556 25050 50820 25060
rect 50652 24612 50708 24622
rect 50652 23716 50708 24556
rect 50652 23660 50932 23716
rect 50556 23548 50820 23558
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50556 23482 50820 23492
rect 50876 23380 50932 23660
rect 50428 23154 50484 23212
rect 50428 23102 50430 23154
rect 50482 23102 50484 23154
rect 50428 23090 50484 23102
rect 50764 23324 50932 23380
rect 50316 22754 50372 22764
rect 49532 22540 49924 22596
rect 49532 22482 49588 22540
rect 49532 22430 49534 22482
rect 49586 22430 49588 22482
rect 49532 22418 49588 22430
rect 50428 22484 50484 22494
rect 49868 22370 49924 22382
rect 49868 22318 49870 22370
rect 49922 22318 49924 22370
rect 49756 22260 49812 22270
rect 49420 22204 49588 22260
rect 49084 21758 49086 21810
rect 49138 21758 49140 21810
rect 49084 21746 49140 21758
rect 49420 21812 49476 21822
rect 49420 21718 49476 21756
rect 48748 21606 48804 21644
rect 48860 21698 48916 21710
rect 48860 21646 48862 21698
rect 48914 21646 48916 21698
rect 48636 21522 48692 21532
rect 48860 20804 48916 21646
rect 49308 21700 49364 21710
rect 49308 21606 49364 21644
rect 49532 21588 49588 22204
rect 49756 22166 49812 22204
rect 49868 21924 49924 22318
rect 50204 22260 50260 22270
rect 50428 22260 50484 22428
rect 50204 22166 50260 22204
rect 50316 22258 50484 22260
rect 50316 22206 50430 22258
rect 50482 22206 50484 22258
rect 50316 22204 50484 22206
rect 49868 21858 49924 21868
rect 49980 22036 50036 22046
rect 49980 21810 50036 21980
rect 49980 21758 49982 21810
rect 50034 21758 50036 21810
rect 49980 21746 50036 21758
rect 48860 20738 48916 20748
rect 49420 21532 49588 21588
rect 49644 21588 49700 21598
rect 49644 21586 49812 21588
rect 49644 21534 49646 21586
rect 49698 21534 49812 21586
rect 49644 21532 49812 21534
rect 49196 20020 49252 20030
rect 48076 19404 48244 19460
rect 48860 20018 49252 20020
rect 48860 19966 49198 20018
rect 49250 19966 49252 20018
rect 48860 19964 49252 19966
rect 47964 19236 48020 19246
rect 47852 19234 48020 19236
rect 47852 19182 47966 19234
rect 48018 19182 48020 19234
rect 47852 19180 48020 19182
rect 48076 19236 48132 19404
rect 48076 19180 48356 19236
rect 47964 19124 48020 19180
rect 47964 19058 48020 19068
rect 48188 19012 48244 19022
rect 48188 18918 48244 18956
rect 47628 17556 47684 17566
rect 47628 16884 47684 17500
rect 48188 17556 48244 17566
rect 48188 17462 48244 17500
rect 48300 17554 48356 19180
rect 48300 17502 48302 17554
rect 48354 17502 48356 17554
rect 48300 17490 48356 17502
rect 48412 19124 48468 19134
rect 48524 19124 48580 19134
rect 48468 19122 48580 19124
rect 48468 19070 48526 19122
rect 48578 19070 48580 19122
rect 48468 19068 48580 19070
rect 47740 17444 47796 17454
rect 47740 17350 47796 17388
rect 47964 17444 48020 17454
rect 47964 17442 48132 17444
rect 47964 17390 47966 17442
rect 48018 17390 48132 17442
rect 47964 17388 48132 17390
rect 47964 17378 48020 17388
rect 47628 15428 47684 16828
rect 47740 16098 47796 16110
rect 47740 16046 47742 16098
rect 47794 16046 47796 16098
rect 47740 15540 47796 16046
rect 48076 16100 48132 17388
rect 48188 16100 48244 16110
rect 48076 16098 48244 16100
rect 48076 16046 48190 16098
rect 48242 16046 48244 16098
rect 48076 16044 48244 16046
rect 48188 16034 48244 16044
rect 47964 15540 48020 15550
rect 47740 15484 47964 15540
rect 47964 15446 48020 15484
rect 47628 15362 47684 15372
rect 47516 15092 47684 15148
rect 46396 14530 46452 15036
rect 46396 14478 46398 14530
rect 46450 14478 46452 14530
rect 46396 14466 46452 14478
rect 46060 14418 46116 14430
rect 46060 14366 46062 14418
rect 46114 14366 46116 14418
rect 46060 14196 46116 14366
rect 46508 14420 46564 14430
rect 46564 14364 46788 14420
rect 46508 14354 46564 14364
rect 46172 14308 46228 14318
rect 46172 14214 46228 14252
rect 46396 14308 46452 14318
rect 46060 14130 46116 14140
rect 46172 13972 46228 13982
rect 45948 12908 46116 12964
rect 45780 12460 45892 12516
rect 45948 12738 46004 12750
rect 45948 12686 45950 12738
rect 46002 12686 46004 12738
rect 45724 12402 45780 12460
rect 45724 12350 45726 12402
rect 45778 12350 45780 12402
rect 45724 12338 45780 12350
rect 45948 11844 46004 12686
rect 45948 11778 46004 11788
rect 45612 11218 45668 11228
rect 45052 10882 45108 10892
rect 45052 10612 45108 10622
rect 45052 10050 45108 10556
rect 45724 10612 45780 10622
rect 45724 10518 45780 10556
rect 45052 9998 45054 10050
rect 45106 9998 45108 10050
rect 45052 9986 45108 9998
rect 45276 10498 45332 10510
rect 45276 10446 45278 10498
rect 45330 10446 45332 10498
rect 45164 9938 45220 9950
rect 45164 9886 45166 9938
rect 45218 9886 45220 9938
rect 45052 9828 45108 9838
rect 45052 9044 45108 9772
rect 45164 9604 45220 9886
rect 45164 9538 45220 9548
rect 45052 8978 45108 8988
rect 45276 8372 45332 10446
rect 45500 10164 45556 10174
rect 45388 9828 45444 9838
rect 45388 9268 45444 9772
rect 45500 9828 45556 10108
rect 46060 10052 46116 12908
rect 46172 12066 46228 13916
rect 46284 12740 46340 12750
rect 46284 12646 46340 12684
rect 46396 12516 46452 14252
rect 46172 12014 46174 12066
rect 46226 12014 46228 12066
rect 46172 11732 46228 12014
rect 46172 11666 46228 11676
rect 46284 12460 46452 12516
rect 46172 10052 46228 10062
rect 46060 9996 46172 10052
rect 46172 9986 46228 9996
rect 45500 9826 45668 9828
rect 45500 9774 45502 9826
rect 45554 9774 45668 9826
rect 45500 9772 45668 9774
rect 45500 9762 45556 9772
rect 45388 9212 45556 9268
rect 45388 9044 45444 9054
rect 45388 8930 45444 8988
rect 45500 9042 45556 9212
rect 45500 8990 45502 9042
rect 45554 8990 45556 9042
rect 45500 8978 45556 8990
rect 45612 9044 45668 9772
rect 46172 9268 46228 9278
rect 46172 9174 46228 9212
rect 45724 9044 45780 9054
rect 45612 9042 45780 9044
rect 45612 8990 45726 9042
rect 45778 8990 45780 9042
rect 45612 8988 45780 8990
rect 45724 8978 45780 8988
rect 45388 8878 45390 8930
rect 45442 8878 45444 8930
rect 45388 8866 45444 8878
rect 45612 8708 45668 8718
rect 45500 8652 45612 8708
rect 45276 8306 45332 8316
rect 45388 8370 45444 8382
rect 45388 8318 45390 8370
rect 45442 8318 45444 8370
rect 45164 8258 45220 8270
rect 45164 8206 45166 8258
rect 45218 8206 45220 8258
rect 45164 7476 45220 8206
rect 45164 6580 45220 7420
rect 45388 8036 45444 8318
rect 45388 6804 45444 7980
rect 45500 7700 45556 8652
rect 45612 8642 45668 8652
rect 45500 7586 45556 7644
rect 45500 7534 45502 7586
rect 45554 7534 45556 7586
rect 45500 7522 45556 7534
rect 45612 8484 45668 8494
rect 45388 6738 45444 6748
rect 45164 6486 45220 6524
rect 45500 6580 45556 6590
rect 45500 6486 45556 6524
rect 44940 6066 44996 6076
rect 45612 5346 45668 8428
rect 45836 8370 45892 8382
rect 45836 8318 45838 8370
rect 45890 8318 45892 8370
rect 45724 7476 45780 7486
rect 45836 7476 45892 8318
rect 45724 7474 45892 7476
rect 45724 7422 45726 7474
rect 45778 7422 45892 7474
rect 45724 7420 45892 7422
rect 46060 7924 46116 7934
rect 46284 7924 46340 12460
rect 46620 11732 46676 11742
rect 46396 10612 46452 10622
rect 46396 10518 46452 10556
rect 46620 10610 46676 11676
rect 46732 10836 46788 14364
rect 46844 14308 46900 14318
rect 46844 14214 46900 14252
rect 46844 13300 46900 13310
rect 46844 13074 46900 13244
rect 46844 13022 46846 13074
rect 46898 13022 46900 13074
rect 46844 13010 46900 13022
rect 46956 12292 47012 15092
rect 46956 12226 47012 12236
rect 47404 13300 47460 13310
rect 46732 10780 47012 10836
rect 46620 10558 46622 10610
rect 46674 10558 46676 10610
rect 46620 10546 46676 10558
rect 46732 10612 46788 10622
rect 46732 10052 46788 10556
rect 46116 7868 46340 7924
rect 46508 9996 46788 10052
rect 45724 7410 45780 7420
rect 46060 6802 46116 7868
rect 46508 7586 46564 9996
rect 46844 9826 46900 9838
rect 46844 9774 46846 9826
rect 46898 9774 46900 9826
rect 46620 9604 46676 9614
rect 46620 9266 46676 9548
rect 46620 9214 46622 9266
rect 46674 9214 46676 9266
rect 46620 9156 46676 9214
rect 46620 9090 46676 9100
rect 46844 8372 46900 9774
rect 46956 9714 47012 10780
rect 47180 10612 47236 10622
rect 47180 10518 47236 10556
rect 46956 9662 46958 9714
rect 47010 9662 47012 9714
rect 46956 9604 47012 9662
rect 46956 9538 47012 9548
rect 47068 10050 47124 10062
rect 47068 9998 47070 10050
rect 47122 9998 47124 10050
rect 46844 8306 46900 8316
rect 47068 7812 47124 9998
rect 47404 9826 47460 13244
rect 47404 9774 47406 9826
rect 47458 9774 47460 9826
rect 47404 9762 47460 9774
rect 47068 7746 47124 7756
rect 46508 7534 46510 7586
rect 46562 7534 46564 7586
rect 46508 7522 46564 7534
rect 46284 7476 46340 7486
rect 46284 7382 46340 7420
rect 46060 6750 46062 6802
rect 46114 6750 46116 6802
rect 46060 6738 46116 6750
rect 46284 6690 46340 6702
rect 46284 6638 46286 6690
rect 46338 6638 46340 6690
rect 45612 5294 45614 5346
rect 45666 5294 45668 5346
rect 45612 5282 45668 5294
rect 46060 6468 46116 6478
rect 44828 5236 44884 5246
rect 44716 5234 44884 5236
rect 44716 5182 44830 5234
rect 44882 5182 44884 5234
rect 44716 5180 44884 5182
rect 44828 5170 44884 5180
rect 46060 5122 46116 6412
rect 46060 5070 46062 5122
rect 46114 5070 46116 5122
rect 46060 5058 46116 5070
rect 46284 5124 46340 6638
rect 46620 6580 46676 6590
rect 46620 5236 46676 6524
rect 46732 6578 46788 6590
rect 46732 6526 46734 6578
rect 46786 6526 46788 6578
rect 46732 6468 46788 6526
rect 47404 6580 47460 6590
rect 47404 6486 47460 6524
rect 46732 6402 46788 6412
rect 47628 5236 47684 15092
rect 48412 11172 48468 19068
rect 48524 19058 48580 19068
rect 48860 19122 48916 19964
rect 49196 19954 49252 19964
rect 49420 19796 49476 21532
rect 49644 21522 49700 21532
rect 49756 20130 49812 21532
rect 50316 21140 50372 22204
rect 50428 22194 50484 22204
rect 50540 22260 50596 22270
rect 50540 22258 50708 22260
rect 50540 22206 50542 22258
rect 50594 22206 50708 22258
rect 50540 22204 50708 22206
rect 50540 22194 50596 22204
rect 50652 22148 50708 22204
rect 50764 22148 50820 23324
rect 50876 23044 50932 23054
rect 50876 22594 50932 22988
rect 50876 22542 50878 22594
rect 50930 22542 50932 22594
rect 50876 22530 50932 22542
rect 51100 23042 51156 23054
rect 51100 22990 51102 23042
rect 51154 22990 51156 23042
rect 51100 22482 51156 22990
rect 51100 22430 51102 22482
rect 51154 22430 51156 22482
rect 51100 22418 51156 22430
rect 51212 22370 51268 25230
rect 51212 22318 51214 22370
rect 51266 22318 51268 22370
rect 50652 22092 50932 22148
rect 50556 21980 50820 21990
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50556 21914 50820 21924
rect 49756 20078 49758 20130
rect 49810 20078 49812 20130
rect 49756 20066 49812 20078
rect 49868 21084 50372 21140
rect 50428 21476 50484 21486
rect 50876 21476 50932 22092
rect 50428 21474 50932 21476
rect 50428 21422 50430 21474
rect 50482 21422 50932 21474
rect 50428 21420 50932 21422
rect 48860 19070 48862 19122
rect 48914 19070 48916 19122
rect 48860 17892 48916 19070
rect 48860 17826 48916 17836
rect 49084 19740 49476 19796
rect 49532 20018 49588 20030
rect 49532 19966 49534 20018
rect 49586 19966 49588 20018
rect 48524 17668 48580 17678
rect 48524 17574 48580 17612
rect 48860 17444 48916 17454
rect 48860 17350 48916 17388
rect 49084 17108 49140 19740
rect 49532 19234 49588 19966
rect 49532 19182 49534 19234
rect 49586 19182 49588 19234
rect 49532 19170 49588 19182
rect 49644 19906 49700 19918
rect 49644 19854 49646 19906
rect 49698 19854 49700 19906
rect 49644 19236 49700 19854
rect 49756 19236 49812 19246
rect 49644 19234 49812 19236
rect 49644 19182 49758 19234
rect 49810 19182 49812 19234
rect 49644 19180 49812 19182
rect 49868 19236 49924 21084
rect 49980 20916 50036 20926
rect 50036 20860 50372 20916
rect 49980 20822 50036 20860
rect 50316 20020 50372 20860
rect 50428 20188 50484 21420
rect 50556 20412 50820 20422
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50556 20346 50820 20356
rect 50428 20132 50596 20188
rect 50428 20020 50484 20030
rect 50316 20018 50484 20020
rect 50316 19966 50430 20018
rect 50482 19966 50484 20018
rect 50316 19964 50484 19966
rect 50204 19908 50260 19918
rect 50092 19852 50204 19908
rect 49980 19236 50036 19246
rect 49868 19234 50036 19236
rect 49868 19182 49982 19234
rect 50034 19182 50036 19234
rect 49868 19180 50036 19182
rect 49756 19170 49812 19180
rect 49980 19170 50036 19180
rect 48972 17052 49140 17108
rect 49196 19122 49252 19134
rect 49196 19070 49198 19122
rect 49250 19070 49252 19122
rect 49196 18452 49252 19070
rect 49308 19010 49364 19022
rect 49308 18958 49310 19010
rect 49362 18958 49364 19010
rect 49308 18900 49364 18958
rect 49308 18834 49364 18844
rect 50092 18900 50148 19852
rect 50204 19842 50260 19852
rect 50204 19124 50260 19134
rect 50204 19030 50260 19068
rect 50316 19122 50372 19134
rect 50316 19070 50318 19122
rect 50370 19070 50372 19122
rect 50316 19012 50372 19070
rect 50316 18946 50372 18956
rect 50092 18562 50148 18844
rect 50428 18676 50484 19964
rect 50540 19796 50596 20132
rect 50540 19730 50596 19740
rect 51100 19906 51156 19918
rect 51100 19854 51102 19906
rect 51154 19854 51156 19906
rect 51100 19458 51156 19854
rect 51100 19406 51102 19458
rect 51154 19406 51156 19458
rect 51100 19394 51156 19406
rect 50988 19236 51044 19246
rect 50764 19124 50820 19134
rect 50764 19030 50820 19068
rect 50988 19124 51044 19180
rect 51212 19124 51268 22318
rect 50988 19122 51268 19124
rect 50988 19070 50990 19122
rect 51042 19070 51268 19122
rect 50988 19068 51268 19070
rect 50988 19058 51044 19068
rect 50556 18844 50820 18854
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50556 18778 50820 18788
rect 50092 18510 50094 18562
rect 50146 18510 50148 18562
rect 50092 18498 50148 18510
rect 50204 18620 50484 18676
rect 50540 18676 50596 18686
rect 49868 18452 49924 18462
rect 49196 17108 49252 18396
rect 49420 18450 49924 18452
rect 49420 18398 49870 18450
rect 49922 18398 49924 18450
rect 49420 18396 49924 18398
rect 49420 17778 49476 18396
rect 49868 18386 49924 18396
rect 49756 17892 49812 17902
rect 49420 17726 49422 17778
rect 49474 17726 49476 17778
rect 49420 17714 49476 17726
rect 49532 17836 49756 17892
rect 49812 17836 49924 17892
rect 49308 17668 49364 17678
rect 49308 17574 49364 17612
rect 48860 16996 48916 17006
rect 48972 16996 49028 17052
rect 49196 17042 49252 17052
rect 48860 16994 49028 16996
rect 48860 16942 48862 16994
rect 48914 16942 49028 16994
rect 48860 16940 49028 16942
rect 48860 16930 48916 16940
rect 48748 16884 48804 16922
rect 48748 16818 48804 16828
rect 49084 16882 49140 16894
rect 49084 16830 49086 16882
rect 49138 16830 49140 16882
rect 49084 16436 49140 16830
rect 49420 16884 49476 16894
rect 49420 16790 49476 16828
rect 49084 16370 49140 16380
rect 48860 16100 48916 16110
rect 49532 16100 49588 17836
rect 49756 17826 49812 17836
rect 49868 17666 49924 17836
rect 49868 17614 49870 17666
rect 49922 17614 49924 17666
rect 49868 17602 49924 17614
rect 49644 17556 49700 17566
rect 49644 17554 49812 17556
rect 49644 17502 49646 17554
rect 49698 17502 49812 17554
rect 49644 17500 49812 17502
rect 49644 17490 49700 17500
rect 49756 17220 49812 17500
rect 49756 17164 50148 17220
rect 49644 17108 49700 17118
rect 49700 17052 49812 17108
rect 49644 17042 49700 17052
rect 49756 16994 49812 17052
rect 50092 17106 50148 17164
rect 50092 17054 50094 17106
rect 50146 17054 50148 17106
rect 50092 17042 50148 17054
rect 49756 16942 49758 16994
rect 49810 16942 49812 16994
rect 49644 16100 49700 16110
rect 48860 16098 49700 16100
rect 48860 16046 48862 16098
rect 48914 16046 49646 16098
rect 49698 16046 49700 16098
rect 48860 16044 49700 16046
rect 48860 16034 48916 16044
rect 49644 16034 49700 16044
rect 48636 15986 48692 15998
rect 48636 15934 48638 15986
rect 48690 15934 48692 15986
rect 48524 15874 48580 15886
rect 48524 15822 48526 15874
rect 48578 15822 48580 15874
rect 48524 14530 48580 15822
rect 48636 15538 48692 15934
rect 49756 15764 49812 16942
rect 49868 16996 49924 17006
rect 49868 16994 50036 16996
rect 49868 16942 49870 16994
rect 49922 16942 50036 16994
rect 49868 16940 50036 16942
rect 49868 16930 49924 16940
rect 49980 16660 50036 16940
rect 50204 16884 50260 18620
rect 50540 18450 50596 18620
rect 51100 18674 51156 19068
rect 51100 18622 51102 18674
rect 51154 18622 51156 18674
rect 51100 18610 51156 18622
rect 50540 18398 50542 18450
rect 50594 18398 50596 18450
rect 50316 18340 50372 18350
rect 50316 18246 50372 18284
rect 50540 17444 50596 18398
rect 50876 18340 50932 18350
rect 50876 18246 50932 18284
rect 51100 18338 51156 18350
rect 51100 18286 51102 18338
rect 51154 18286 51156 18338
rect 50540 17388 50932 17444
rect 50556 17276 50820 17286
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50556 17210 50820 17220
rect 50316 16884 50372 16894
rect 50260 16882 50372 16884
rect 50260 16830 50318 16882
rect 50370 16830 50372 16882
rect 50260 16828 50372 16830
rect 50204 16790 50260 16828
rect 49980 16594 50036 16604
rect 49980 16436 50036 16446
rect 50036 16380 50260 16436
rect 49980 16370 50036 16380
rect 49980 16212 50036 16222
rect 48636 15486 48638 15538
rect 48690 15486 48692 15538
rect 48636 15474 48692 15486
rect 49532 15708 49812 15764
rect 49868 15986 49924 15998
rect 49868 15934 49870 15986
rect 49922 15934 49924 15986
rect 48860 15428 48916 15438
rect 48748 15426 48916 15428
rect 48748 15374 48862 15426
rect 48914 15374 48916 15426
rect 48748 15372 48916 15374
rect 48748 15092 48804 15372
rect 48860 15362 48916 15372
rect 48972 15428 49028 15438
rect 49532 15428 49588 15708
rect 49868 15538 49924 15934
rect 49868 15486 49870 15538
rect 49922 15486 49924 15538
rect 49868 15474 49924 15486
rect 48972 15426 49588 15428
rect 48972 15374 48974 15426
rect 49026 15374 49534 15426
rect 49586 15374 49588 15426
rect 48972 15372 49588 15374
rect 48972 15362 49028 15372
rect 49532 15362 49588 15372
rect 49644 15426 49700 15438
rect 49644 15374 49646 15426
rect 49698 15374 49700 15426
rect 48524 14478 48526 14530
rect 48578 14478 48580 14530
rect 48524 14466 48580 14478
rect 48636 15036 48804 15092
rect 49084 15092 49140 15102
rect 48636 13300 48692 15036
rect 48860 14532 48916 14570
rect 48860 14466 48916 14476
rect 49084 14530 49140 15036
rect 49084 14478 49086 14530
rect 49138 14478 49140 14530
rect 49084 14466 49140 14478
rect 49644 14532 49700 15374
rect 49980 14644 50036 16156
rect 50204 16098 50260 16380
rect 50204 16046 50206 16098
rect 50258 16046 50260 16098
rect 50204 16034 50260 16046
rect 50092 15874 50148 15886
rect 50092 15822 50094 15874
rect 50146 15822 50148 15874
rect 50092 15426 50148 15822
rect 50316 15764 50372 16828
rect 50092 15374 50094 15426
rect 50146 15374 50148 15426
rect 50092 15362 50148 15374
rect 50204 15708 50372 15764
rect 50556 15708 50820 15718
rect 50204 15540 50260 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50556 15642 50820 15652
rect 49980 14578 50036 14588
rect 48636 13234 48692 13244
rect 48860 14306 48916 14318
rect 48860 14254 48862 14306
rect 48914 14254 48916 14306
rect 48860 13076 48916 14254
rect 48748 13020 48916 13076
rect 49084 14308 49140 14318
rect 48748 12290 48804 13020
rect 48972 12852 49028 12862
rect 48860 12850 49028 12852
rect 48860 12798 48974 12850
rect 49026 12798 49028 12850
rect 48860 12796 49028 12798
rect 48860 12402 48916 12796
rect 48972 12786 49028 12796
rect 48860 12350 48862 12402
rect 48914 12350 48916 12402
rect 48860 12338 48916 12350
rect 48972 12516 49028 12526
rect 48748 12238 48750 12290
rect 48802 12238 48804 12290
rect 48748 12226 48804 12238
rect 48972 12290 49028 12460
rect 48972 12238 48974 12290
rect 49026 12238 49028 12290
rect 48972 11844 49028 12238
rect 48972 11778 49028 11788
rect 48860 11284 48916 11294
rect 49084 11284 49140 14252
rect 49644 13636 49700 14476
rect 49644 13570 49700 13580
rect 49980 13636 50036 13646
rect 50204 13636 50260 15484
rect 50428 15538 50484 15550
rect 50428 15486 50430 15538
rect 50482 15486 50484 15538
rect 50316 15316 50372 15326
rect 50316 15222 50372 15260
rect 50316 13746 50372 13758
rect 50316 13694 50318 13746
rect 50370 13694 50372 13746
rect 50316 13636 50372 13694
rect 49980 13634 50372 13636
rect 49980 13582 49982 13634
rect 50034 13582 50372 13634
rect 49980 13580 50372 13582
rect 49756 12962 49812 12974
rect 49756 12910 49758 12962
rect 49810 12910 49812 12962
rect 49756 12740 49812 12910
rect 49980 12740 50036 13580
rect 50428 13188 50484 15486
rect 50652 15316 50708 15326
rect 50876 15316 50932 17388
rect 51100 16994 51156 18286
rect 52332 17444 52388 29932
rect 52892 29922 52948 29932
rect 53116 29316 53172 31724
rect 53228 31556 53284 31566
rect 53228 30882 53284 31500
rect 53228 30830 53230 30882
rect 53282 30830 53284 30882
rect 53228 30818 53284 30830
rect 53228 30100 53284 30110
rect 53228 30006 53284 30044
rect 53228 29316 53284 29326
rect 53116 29314 53284 29316
rect 53116 29262 53230 29314
rect 53282 29262 53284 29314
rect 53116 29260 53284 29262
rect 53228 29250 53284 29260
rect 52892 27970 52948 27982
rect 52892 27918 52894 27970
rect 52946 27918 52948 27970
rect 52668 27746 52724 27758
rect 52668 27694 52670 27746
rect 52722 27694 52724 27746
rect 52668 27412 52724 27694
rect 52668 27346 52724 27356
rect 52892 26908 52948 27918
rect 53228 27858 53284 27870
rect 53228 27806 53230 27858
rect 53282 27806 53284 27858
rect 53228 27412 53284 27806
rect 53228 27346 53284 27356
rect 52556 26852 52948 26908
rect 52556 24052 52612 26852
rect 53228 26178 53284 26190
rect 53228 26126 53230 26178
rect 53282 26126 53284 26178
rect 53228 25620 53284 26126
rect 53228 25554 53284 25564
rect 53228 25394 53284 25406
rect 53228 25342 53230 25394
rect 53282 25342 53284 25394
rect 52556 23986 52612 23996
rect 52892 25282 52948 25294
rect 52892 25230 52894 25282
rect 52946 25230 52948 25282
rect 52892 23940 52948 25230
rect 53228 24724 53284 25342
rect 53228 24630 53284 24668
rect 52892 23874 52948 23884
rect 53228 23042 53284 23054
rect 53228 22990 53230 23042
rect 53282 22990 53284 23042
rect 53228 22484 53284 22990
rect 53228 22418 53284 22428
rect 53228 22258 53284 22270
rect 53228 22206 53230 22258
rect 53282 22206 53284 22258
rect 52892 22146 52948 22158
rect 52892 22094 52894 22146
rect 52946 22094 52948 22146
rect 52892 21812 52948 22094
rect 53228 22036 53284 22206
rect 53340 22036 53396 22046
rect 53228 21980 53340 22036
rect 52892 21746 52948 21756
rect 53340 21810 53396 21980
rect 53340 21758 53342 21810
rect 53394 21758 53396 21810
rect 53340 21746 53396 21758
rect 52332 17378 52388 17388
rect 52780 21588 52836 21598
rect 51100 16942 51102 16994
rect 51154 16942 51156 16994
rect 51100 16930 51156 16942
rect 50652 15314 50932 15316
rect 50652 15262 50654 15314
rect 50706 15262 50932 15314
rect 50652 15260 50932 15262
rect 50988 16772 51044 16782
rect 50988 15316 51044 16716
rect 52780 15988 52836 21532
rect 52892 20804 52948 20814
rect 52892 19122 52948 20748
rect 53228 19908 53284 19918
rect 53228 19814 53284 19852
rect 52892 19070 52894 19122
rect 52946 19070 52948 19122
rect 52892 19058 52948 19070
rect 53228 19348 53284 19358
rect 53228 19234 53284 19292
rect 53228 19182 53230 19234
rect 53282 19182 53284 19234
rect 53228 18676 53284 19182
rect 53340 18676 53396 18686
rect 53228 18674 53396 18676
rect 53228 18622 53342 18674
rect 53394 18622 53396 18674
rect 53228 18620 53396 18622
rect 53340 18610 53396 18620
rect 53228 16772 53284 16782
rect 53228 16678 53284 16716
rect 53116 16660 53172 16670
rect 53116 16100 53172 16604
rect 53116 16098 53396 16100
rect 53116 16046 53118 16098
rect 53170 16046 53396 16098
rect 53116 16044 53396 16046
rect 53116 16034 53172 16044
rect 52892 15988 52948 15998
rect 52780 15986 52948 15988
rect 52780 15934 52894 15986
rect 52946 15934 52948 15986
rect 52780 15932 52948 15934
rect 52892 15922 52948 15932
rect 53340 15538 53396 16044
rect 53340 15486 53342 15538
rect 53394 15486 53396 15538
rect 53340 15474 53396 15486
rect 50652 15204 50708 15260
rect 50988 15250 51044 15260
rect 50652 15138 50708 15148
rect 52668 14644 52724 14654
rect 52668 14550 52724 14588
rect 52220 14306 52276 14318
rect 52220 14254 52222 14306
rect 52274 14254 52276 14306
rect 50556 14140 50820 14150
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50556 14074 50820 14084
rect 52220 13972 52276 14254
rect 52220 13906 52276 13916
rect 53228 14306 53284 14318
rect 53228 14254 53230 14306
rect 53282 14254 53284 14306
rect 53228 13972 53284 14254
rect 53228 13906 53284 13916
rect 51100 13636 51156 13646
rect 50876 13634 51156 13636
rect 50876 13582 51102 13634
rect 51154 13582 51156 13634
rect 50876 13580 51156 13582
rect 50540 13188 50596 13198
rect 50428 13186 50596 13188
rect 50428 13134 50542 13186
rect 50594 13134 50596 13186
rect 50428 13132 50596 13134
rect 50540 13122 50596 13132
rect 50876 13186 50932 13580
rect 51100 13570 51156 13580
rect 53228 13636 53284 13646
rect 53228 13542 53284 13580
rect 50876 13134 50878 13186
rect 50930 13134 50932 13186
rect 50876 13122 50932 13134
rect 50204 12740 50260 12750
rect 49756 12738 50260 12740
rect 49756 12686 50206 12738
rect 50258 12686 50260 12738
rect 49756 12684 50260 12686
rect 48860 11282 49700 11284
rect 48860 11230 48862 11282
rect 48914 11230 49700 11282
rect 48860 11228 49700 11230
rect 48860 11218 48916 11228
rect 48524 11172 48580 11182
rect 48412 11170 48580 11172
rect 48412 11118 48526 11170
rect 48578 11118 48580 11170
rect 48412 11116 48580 11118
rect 47964 9826 48020 9838
rect 47964 9774 47966 9826
rect 48018 9774 48020 9826
rect 47964 9716 48020 9774
rect 47964 9650 48020 9660
rect 48524 9268 48580 11116
rect 48972 10780 49588 10836
rect 48972 10498 49028 10780
rect 49196 10612 49252 10622
rect 48972 10446 48974 10498
rect 49026 10446 49028 10498
rect 48860 9828 48916 9838
rect 48860 9714 48916 9772
rect 48860 9662 48862 9714
rect 48914 9662 48916 9714
rect 48860 9650 48916 9662
rect 48524 9202 48580 9212
rect 48748 8930 48804 8942
rect 48748 8878 48750 8930
rect 48802 8878 48804 8930
rect 48636 8372 48692 8382
rect 47740 8260 47796 8270
rect 47740 8166 47796 8204
rect 48076 8146 48132 8158
rect 48076 8094 48078 8146
rect 48130 8094 48132 8146
rect 48076 7698 48132 8094
rect 48636 8148 48692 8316
rect 48748 8260 48804 8878
rect 48860 8260 48916 8270
rect 48748 8258 48916 8260
rect 48748 8206 48862 8258
rect 48914 8206 48916 8258
rect 48748 8204 48916 8206
rect 48860 8194 48916 8204
rect 48972 8260 49028 10446
rect 49084 10556 49196 10612
rect 49084 8708 49140 10556
rect 49196 10518 49252 10556
rect 49420 10610 49476 10622
rect 49420 10558 49422 10610
rect 49474 10558 49476 10610
rect 49308 10498 49364 10510
rect 49308 10446 49310 10498
rect 49362 10446 49364 10498
rect 49308 9940 49364 10446
rect 49308 9874 49364 9884
rect 49420 9940 49476 10558
rect 49532 10388 49588 10780
rect 49644 10610 49700 11228
rect 49980 11170 50036 11182
rect 49980 11118 49982 11170
rect 50034 11118 50036 11170
rect 49644 10558 49646 10610
rect 49698 10558 49700 10610
rect 49644 10546 49700 10558
rect 49756 10610 49812 10622
rect 49756 10558 49758 10610
rect 49810 10558 49812 10610
rect 49756 10388 49812 10558
rect 49980 10612 50036 11118
rect 50204 10612 50260 12684
rect 50764 12740 50820 12778
rect 50764 12674 50820 12684
rect 50556 12572 50820 12582
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50556 12506 50820 12516
rect 52444 12292 52500 12302
rect 52444 12198 52500 12236
rect 52780 12068 52836 12078
rect 52780 12066 52948 12068
rect 52780 12014 52782 12066
rect 52834 12014 52948 12066
rect 52780 12012 52948 12014
rect 52780 12002 52836 12012
rect 52892 11282 52948 12012
rect 53340 12066 53396 12078
rect 53340 12014 53342 12066
rect 53394 12014 53396 12066
rect 52892 11230 52894 11282
rect 52946 11230 52948 11282
rect 52892 11218 52948 11230
rect 53228 11284 53284 11294
rect 53340 11284 53396 12014
rect 53284 11228 53396 11284
rect 53228 11190 53284 11228
rect 50556 11004 50820 11014
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50556 10938 50820 10948
rect 50316 10612 50372 10622
rect 49980 10610 50372 10612
rect 49980 10558 50318 10610
rect 50370 10558 50372 10610
rect 49980 10556 50372 10558
rect 49532 10332 49812 10388
rect 49420 9884 49812 9940
rect 49420 9828 49476 9884
rect 49420 9762 49476 9772
rect 49196 9716 49252 9726
rect 49196 9622 49252 9660
rect 49532 9714 49588 9726
rect 49532 9662 49534 9714
rect 49586 9662 49588 9714
rect 49532 9604 49588 9662
rect 49420 9548 49532 9604
rect 49420 9042 49476 9548
rect 49532 9538 49588 9548
rect 49420 8990 49422 9042
rect 49474 8990 49476 9042
rect 49420 8978 49476 8990
rect 49532 8930 49588 8942
rect 49532 8878 49534 8930
rect 49586 8878 49588 8930
rect 49084 8652 49364 8708
rect 49084 8260 49140 8270
rect 48972 8204 49084 8260
rect 48636 8146 48804 8148
rect 48636 8094 48638 8146
rect 48690 8094 48804 8146
rect 48636 8092 48804 8094
rect 48636 8082 48692 8092
rect 48188 8036 48244 8046
rect 48188 7942 48244 7980
rect 48412 8034 48468 8046
rect 48412 7982 48414 8034
rect 48466 7982 48468 8034
rect 48076 7646 48078 7698
rect 48130 7646 48132 7698
rect 48076 7634 48132 7646
rect 47740 7586 47796 7598
rect 47740 7534 47742 7586
rect 47794 7534 47796 7586
rect 47740 6804 47796 7534
rect 47964 7588 48020 7598
rect 47964 7494 48020 7532
rect 48188 7476 48244 7486
rect 48188 7382 48244 7420
rect 47740 6738 47796 6748
rect 48188 6804 48244 6814
rect 46620 5234 47124 5236
rect 46620 5182 46622 5234
rect 46674 5182 47124 5234
rect 46620 5180 47124 5182
rect 46620 5170 46676 5180
rect 46284 5030 46340 5068
rect 46508 5124 46564 5134
rect 46508 5010 46564 5068
rect 46508 4958 46510 5010
rect 46562 4958 46564 5010
rect 46508 4946 46564 4958
rect 44940 4898 44996 4910
rect 44940 4846 44942 4898
rect 44994 4846 44996 4898
rect 44940 4450 44996 4846
rect 44940 4398 44942 4450
rect 44994 4398 44996 4450
rect 44940 4386 44996 4398
rect 44268 4340 44324 4350
rect 44268 4246 44324 4284
rect 47068 4226 47124 5180
rect 47628 5234 47908 5236
rect 47628 5182 47630 5234
rect 47682 5182 47908 5234
rect 47628 5180 47908 5182
rect 47628 5170 47684 5180
rect 47852 4450 47908 5180
rect 48188 5234 48244 6748
rect 48412 6692 48468 7982
rect 48524 8036 48580 8046
rect 48524 7700 48580 7980
rect 48636 7700 48692 7710
rect 48524 7698 48692 7700
rect 48524 7646 48638 7698
rect 48690 7646 48692 7698
rect 48524 7644 48692 7646
rect 48636 7634 48692 7644
rect 48748 7028 48804 8092
rect 48748 6962 48804 6972
rect 48412 6626 48468 6636
rect 48972 6916 49028 8204
rect 49084 8166 49140 8204
rect 48972 6356 49028 6860
rect 49084 7250 49140 7262
rect 49084 7198 49086 7250
rect 49138 7198 49140 7250
rect 49084 6804 49140 7198
rect 49196 7252 49252 8652
rect 49308 8370 49364 8652
rect 49308 8318 49310 8370
rect 49362 8318 49364 8370
rect 49308 8306 49364 8318
rect 49532 8148 49588 8878
rect 49420 8146 49588 8148
rect 49420 8094 49534 8146
rect 49586 8094 49588 8146
rect 49420 8092 49588 8094
rect 49420 7812 49476 8092
rect 49532 8082 49588 8092
rect 49644 8036 49700 8046
rect 49644 7942 49700 7980
rect 49308 7476 49364 7486
rect 49420 7476 49476 7756
rect 49364 7420 49476 7476
rect 49532 7588 49588 7598
rect 49532 7476 49588 7532
rect 49756 7476 49812 9884
rect 49868 9716 49924 9726
rect 49868 9622 49924 9660
rect 49532 7474 49812 7476
rect 49532 7422 49534 7474
rect 49586 7422 49812 7474
rect 49532 7420 49812 7422
rect 49980 7476 50036 7486
rect 50316 7476 50372 10556
rect 51100 10500 51156 10510
rect 50876 10498 51156 10500
rect 50876 10446 51102 10498
rect 51154 10446 51156 10498
rect 50876 10444 51156 10446
rect 50876 10050 50932 10444
rect 51100 10434 51156 10444
rect 53228 10500 53284 10510
rect 53228 10498 53396 10500
rect 53228 10446 53230 10498
rect 53282 10446 53396 10498
rect 53228 10444 53396 10446
rect 53228 10434 53284 10444
rect 50876 9998 50878 10050
rect 50930 9998 50932 10050
rect 50876 9986 50932 9998
rect 52892 10052 52948 10062
rect 50764 9940 50820 9950
rect 50764 9846 50820 9884
rect 50556 9436 50820 9446
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50556 9370 50820 9380
rect 52892 9266 52948 9996
rect 52892 9214 52894 9266
rect 52946 9214 52948 9266
rect 52892 9202 52948 9214
rect 53340 9716 53396 10444
rect 53228 9042 53284 9054
rect 53228 8990 53230 9042
rect 53282 8990 53284 9042
rect 52668 8932 52724 8942
rect 53228 8932 53284 8990
rect 52668 8930 53284 8932
rect 52668 8878 52670 8930
rect 52722 8878 53284 8930
rect 52668 8876 53284 8878
rect 52668 8866 52724 8876
rect 53228 8596 53284 8876
rect 53228 8530 53284 8540
rect 50540 8148 50596 8158
rect 50540 8054 50596 8092
rect 50652 8036 50708 8046
rect 52668 8036 52724 8046
rect 50652 8034 51156 8036
rect 50652 7982 50654 8034
rect 50706 7982 51156 8034
rect 50652 7980 51156 7982
rect 50652 7970 50708 7980
rect 50556 7868 50820 7878
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50556 7802 50820 7812
rect 51100 7586 51156 7980
rect 52668 7942 52724 7980
rect 53004 8036 53060 8046
rect 53004 8034 53284 8036
rect 53004 7982 53006 8034
rect 53058 7982 53284 8034
rect 53004 7980 53284 7982
rect 51100 7534 51102 7586
rect 51154 7534 51156 7586
rect 51100 7522 51156 7534
rect 49980 7474 50372 7476
rect 49980 7422 49982 7474
rect 50034 7422 50318 7474
rect 50370 7422 50372 7474
rect 49980 7420 50372 7422
rect 49308 7382 49364 7420
rect 49532 7410 49588 7420
rect 49980 7410 50036 7420
rect 49196 7196 50148 7252
rect 49084 6690 49140 6748
rect 49084 6638 49086 6690
rect 49138 6638 49140 6690
rect 49084 6626 49140 6638
rect 49308 7028 49364 7038
rect 49308 6690 49364 6972
rect 49868 6916 49924 6926
rect 49868 6822 49924 6860
rect 50092 6802 50148 7196
rect 50092 6750 50094 6802
rect 50146 6750 50148 6802
rect 50092 6738 50148 6750
rect 49308 6638 49310 6690
rect 49362 6638 49364 6690
rect 49308 6626 49364 6638
rect 49644 6692 49700 6702
rect 49644 6598 49700 6636
rect 49868 6466 49924 6478
rect 49868 6414 49870 6466
rect 49922 6414 49924 6466
rect 48972 6300 49252 6356
rect 49196 6130 49252 6300
rect 49196 6078 49198 6130
rect 49250 6078 49252 6130
rect 49196 6066 49252 6078
rect 49868 6018 49924 6414
rect 49868 5966 49870 6018
rect 49922 5966 49924 6018
rect 49868 5954 49924 5966
rect 50204 5908 50260 7420
rect 50316 7410 50372 7420
rect 53004 6914 53060 7980
rect 53228 7362 53284 7980
rect 53228 7310 53230 7362
rect 53282 7310 53284 7362
rect 53228 7298 53284 7310
rect 53004 6862 53006 6914
rect 53058 6862 53060 6914
rect 53004 6850 53060 6862
rect 50316 6804 50372 6814
rect 50316 6690 50372 6748
rect 53228 6804 53284 6814
rect 53340 6804 53396 9660
rect 53228 6802 53396 6804
rect 53228 6750 53230 6802
rect 53282 6750 53396 6802
rect 53228 6748 53396 6750
rect 53228 6738 53284 6748
rect 50316 6638 50318 6690
rect 50370 6638 50372 6690
rect 50316 6626 50372 6638
rect 51548 6690 51604 6702
rect 51548 6638 51550 6690
rect 51602 6638 51604 6690
rect 51324 6468 51380 6478
rect 51324 6374 51380 6412
rect 50556 6300 50820 6310
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50556 6234 50820 6244
rect 51548 6132 51604 6638
rect 51548 6066 51604 6076
rect 51996 6690 52052 6702
rect 51996 6638 51998 6690
rect 52050 6638 52052 6690
rect 51996 6468 52052 6638
rect 52668 6580 52724 6590
rect 52668 6486 52724 6524
rect 50316 5908 50372 5918
rect 50204 5906 50372 5908
rect 50204 5854 50318 5906
rect 50370 5854 50372 5906
rect 50204 5852 50372 5854
rect 48188 5182 48190 5234
rect 48242 5182 48244 5234
rect 48188 5170 48244 5182
rect 49532 5794 49588 5806
rect 49532 5742 49534 5794
rect 49586 5742 49588 5794
rect 48636 5124 48692 5134
rect 48636 5030 48692 5068
rect 49084 5124 49140 5134
rect 49532 5124 49588 5742
rect 49980 5684 50036 5694
rect 49980 5590 50036 5628
rect 49084 5122 49588 5124
rect 49084 5070 49086 5122
rect 49138 5070 49588 5122
rect 49084 5068 49588 5070
rect 47852 4398 47854 4450
rect 47906 4398 47908 4450
rect 47852 4386 47908 4398
rect 48188 4452 48244 4462
rect 48188 4358 48244 4396
rect 47516 4340 47572 4350
rect 47516 4246 47572 4284
rect 49084 4340 49140 5068
rect 49084 4274 49140 4284
rect 50316 4340 50372 5852
rect 51996 5908 52052 6412
rect 51996 5842 52052 5852
rect 51100 5796 51156 5806
rect 51100 5702 51156 5740
rect 53228 5794 53284 5806
rect 53228 5742 53230 5794
rect 53282 5742 53284 5794
rect 53228 5124 53284 5742
rect 53228 5058 53284 5068
rect 52668 5012 52724 5022
rect 50556 4732 50820 4742
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50556 4666 50820 4676
rect 50876 4452 50932 4462
rect 50876 4358 50932 4396
rect 50316 4274 50372 4284
rect 51660 4340 51716 4350
rect 51660 4246 51716 4284
rect 47068 4174 47070 4226
rect 47122 4174 47124 4226
rect 47068 4162 47124 4174
rect 48748 4226 48804 4238
rect 48748 4174 48750 4226
rect 48802 4174 48804 4226
rect 46956 3556 47012 3566
rect 46956 3462 47012 3500
rect 47628 3556 47684 3566
rect 43932 3442 44212 3444
rect 43932 3390 43934 3442
rect 43986 3390 44212 3442
rect 43932 3388 44212 3390
rect 47628 3388 47684 3500
rect 48524 3556 48580 3566
rect 48748 3556 48804 4174
rect 50428 3668 50484 3678
rect 50428 3574 50484 3612
rect 51996 3668 52052 3678
rect 48524 3554 48804 3556
rect 48524 3502 48526 3554
rect 48578 3502 48804 3554
rect 48524 3500 48804 3502
rect 48524 3490 48580 3500
rect 43932 3378 43988 3388
rect 47404 3332 47460 3342
rect 47404 3238 47460 3276
rect 47516 3332 47684 3388
rect 47516 800 47572 3332
rect 50556 3164 50820 3174
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50556 3098 50820 3108
rect 51996 800 52052 3612
rect 52668 3666 52724 4956
rect 52668 3614 52670 3666
rect 52722 3614 52724 3666
rect 52668 3602 52724 3614
rect 52444 3442 52500 3454
rect 52444 3390 52446 3442
rect 52498 3390 52500 3442
rect 52444 3220 52500 3390
rect 52444 3154 52500 3164
rect 53228 3442 53284 3454
rect 53228 3390 53230 3442
rect 53282 3390 53284 3442
rect 53228 3220 53284 3390
rect 53228 3154 53284 3164
rect 2688 0 2800 800
rect 7168 0 7280 800
rect 11648 0 11760 800
rect 16128 0 16240 800
rect 20608 0 20720 800
rect 25088 0 25200 800
rect 29568 0 29680 800
rect 34048 0 34160 800
rect 38528 0 38640 800
rect 43008 0 43120 800
rect 47488 0 47600 800
rect 51968 0 52080 800
<< via2 >>
rect 4476 50986 4532 50988
rect 4476 50934 4478 50986
rect 4478 50934 4530 50986
rect 4530 50934 4532 50986
rect 4476 50932 4532 50934
rect 4580 50986 4636 50988
rect 4580 50934 4582 50986
rect 4582 50934 4634 50986
rect 4634 50934 4636 50986
rect 4580 50932 4636 50934
rect 4684 50986 4740 50988
rect 4684 50934 4686 50986
rect 4686 50934 4738 50986
rect 4738 50934 4740 50986
rect 4684 50932 4740 50934
rect 19836 51770 19892 51772
rect 19836 51718 19838 51770
rect 19838 51718 19890 51770
rect 19890 51718 19892 51770
rect 19836 51716 19892 51718
rect 19940 51770 19996 51772
rect 19940 51718 19942 51770
rect 19942 51718 19994 51770
rect 19994 51718 19996 51770
rect 19940 51716 19996 51718
rect 20044 51770 20100 51772
rect 20044 51718 20046 51770
rect 20046 51718 20098 51770
rect 20098 51718 20100 51770
rect 20044 51716 20100 51718
rect 50556 51770 50612 51772
rect 50556 51718 50558 51770
rect 50558 51718 50610 51770
rect 50610 51718 50612 51770
rect 50556 51716 50612 51718
rect 50660 51770 50716 51772
rect 50660 51718 50662 51770
rect 50662 51718 50714 51770
rect 50714 51718 50716 51770
rect 50660 51716 50716 51718
rect 50764 51770 50820 51772
rect 50764 51718 50766 51770
rect 50766 51718 50818 51770
rect 50818 51718 50820 51770
rect 50764 51716 50820 51718
rect 51100 51548 51156 51604
rect 35196 50986 35252 50988
rect 35196 50934 35198 50986
rect 35198 50934 35250 50986
rect 35250 50934 35252 50986
rect 35196 50932 35252 50934
rect 35300 50986 35356 50988
rect 35300 50934 35302 50986
rect 35302 50934 35354 50986
rect 35354 50934 35356 50986
rect 35300 50932 35356 50934
rect 35404 50986 35460 50988
rect 35404 50934 35406 50986
rect 35406 50934 35458 50986
rect 35458 50934 35460 50986
rect 35404 50932 35460 50934
rect 49644 51324 49700 51380
rect 13692 50316 13748 50372
rect 13580 49644 13636 49700
rect 4476 49418 4532 49420
rect 4476 49366 4478 49418
rect 4478 49366 4530 49418
rect 4530 49366 4532 49418
rect 4476 49364 4532 49366
rect 4580 49418 4636 49420
rect 4580 49366 4582 49418
rect 4582 49366 4634 49418
rect 4634 49366 4636 49418
rect 4580 49364 4636 49366
rect 4684 49418 4740 49420
rect 4684 49366 4686 49418
rect 4686 49366 4738 49418
rect 4738 49366 4740 49418
rect 4684 49364 4740 49366
rect 16380 50482 16436 50484
rect 16380 50430 16382 50482
rect 16382 50430 16434 50482
rect 16434 50430 16436 50482
rect 16380 50428 16436 50430
rect 17724 50428 17780 50484
rect 20748 50428 20804 50484
rect 15708 49644 15764 49700
rect 16492 49644 16548 49700
rect 4476 47850 4532 47852
rect 4476 47798 4478 47850
rect 4478 47798 4530 47850
rect 4530 47798 4532 47850
rect 4476 47796 4532 47798
rect 4580 47850 4636 47852
rect 4580 47798 4582 47850
rect 4582 47798 4634 47850
rect 4634 47798 4636 47850
rect 4580 47796 4636 47798
rect 4684 47850 4740 47852
rect 4684 47798 4686 47850
rect 4686 47798 4738 47850
rect 4738 47798 4740 47850
rect 4684 47796 4740 47798
rect 11340 47404 11396 47460
rect 4476 46282 4532 46284
rect 4476 46230 4478 46282
rect 4478 46230 4530 46282
rect 4530 46230 4532 46282
rect 4476 46228 4532 46230
rect 4580 46282 4636 46284
rect 4580 46230 4582 46282
rect 4582 46230 4634 46282
rect 4634 46230 4636 46282
rect 4580 46228 4636 46230
rect 4684 46282 4740 46284
rect 4684 46230 4686 46282
rect 4686 46230 4738 46282
rect 4738 46230 4740 46282
rect 4684 46228 4740 46230
rect 4476 44714 4532 44716
rect 4476 44662 4478 44714
rect 4478 44662 4530 44714
rect 4530 44662 4532 44714
rect 4476 44660 4532 44662
rect 4580 44714 4636 44716
rect 4580 44662 4582 44714
rect 4582 44662 4634 44714
rect 4634 44662 4636 44714
rect 4580 44660 4636 44662
rect 4684 44714 4740 44716
rect 4684 44662 4686 44714
rect 4686 44662 4738 44714
rect 4738 44662 4740 44714
rect 4684 44660 4740 44662
rect 4476 43146 4532 43148
rect 4476 43094 4478 43146
rect 4478 43094 4530 43146
rect 4530 43094 4532 43146
rect 4476 43092 4532 43094
rect 4580 43146 4636 43148
rect 4580 43094 4582 43146
rect 4582 43094 4634 43146
rect 4634 43094 4636 43146
rect 4580 43092 4636 43094
rect 4684 43146 4740 43148
rect 4684 43094 4686 43146
rect 4686 43094 4738 43146
rect 4738 43094 4740 43146
rect 4684 43092 4740 43094
rect 9436 45276 9492 45332
rect 14028 47458 14084 47460
rect 14028 47406 14030 47458
rect 14030 47406 14082 47458
rect 14082 47406 14084 47458
rect 14028 47404 14084 47406
rect 13244 47292 13300 47348
rect 14140 47346 14196 47348
rect 14140 47294 14142 47346
rect 14142 47294 14194 47346
rect 14194 47294 14196 47346
rect 14140 47292 14196 47294
rect 11564 45500 11620 45556
rect 11564 45330 11620 45332
rect 11564 45278 11566 45330
rect 11566 45278 11618 45330
rect 11618 45278 11620 45330
rect 11564 45276 11620 45278
rect 12236 46786 12292 46788
rect 12236 46734 12238 46786
rect 12238 46734 12290 46786
rect 12290 46734 12292 46786
rect 12236 46732 12292 46734
rect 14028 46786 14084 46788
rect 14028 46734 14030 46786
rect 14030 46734 14082 46786
rect 14082 46734 14084 46786
rect 14028 46732 14084 46734
rect 12348 46674 12404 46676
rect 12348 46622 12350 46674
rect 12350 46622 12402 46674
rect 12402 46622 12404 46674
rect 12348 46620 12404 46622
rect 11788 45218 11844 45220
rect 11788 45166 11790 45218
rect 11790 45166 11842 45218
rect 11842 45166 11844 45218
rect 11788 45164 11844 45166
rect 10892 43538 10948 43540
rect 10892 43486 10894 43538
rect 10894 43486 10946 43538
rect 10946 43486 10948 43538
rect 10892 43484 10948 43486
rect 9660 43372 9716 43428
rect 5068 41804 5124 41860
rect 4476 41578 4532 41580
rect 4476 41526 4478 41578
rect 4478 41526 4530 41578
rect 4530 41526 4532 41578
rect 4476 41524 4532 41526
rect 4580 41578 4636 41580
rect 4580 41526 4582 41578
rect 4582 41526 4634 41578
rect 4634 41526 4636 41578
rect 4580 41524 4636 41526
rect 4684 41578 4740 41580
rect 4684 41526 4686 41578
rect 4686 41526 4738 41578
rect 4738 41526 4740 41578
rect 4684 41524 4740 41526
rect 4476 40010 4532 40012
rect 4476 39958 4478 40010
rect 4478 39958 4530 40010
rect 4530 39958 4532 40010
rect 4476 39956 4532 39958
rect 4580 40010 4636 40012
rect 4580 39958 4582 40010
rect 4582 39958 4634 40010
rect 4634 39958 4636 40010
rect 4580 39956 4636 39958
rect 4684 40010 4740 40012
rect 4684 39958 4686 40010
rect 4686 39958 4738 40010
rect 4738 39958 4740 40010
rect 4684 39956 4740 39958
rect 8316 41858 8372 41860
rect 8316 41806 8318 41858
rect 8318 41806 8370 41858
rect 8370 41806 8372 41858
rect 8316 41804 8372 41806
rect 8876 41804 8932 41860
rect 9884 41804 9940 41860
rect 5068 39676 5124 39732
rect 4956 39506 5012 39508
rect 4956 39454 4958 39506
rect 4958 39454 5010 39506
rect 5010 39454 5012 39506
rect 4956 39452 5012 39454
rect 5068 39394 5124 39396
rect 5068 39342 5070 39394
rect 5070 39342 5122 39394
rect 5122 39342 5124 39394
rect 5068 39340 5124 39342
rect 5516 39340 5572 39396
rect 6076 39340 6132 39396
rect 5404 38556 5460 38612
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 2492 37154 2548 37156
rect 2492 37102 2494 37154
rect 2494 37102 2546 37154
rect 2546 37102 2548 37154
rect 2492 37100 2548 37102
rect 5068 37772 5124 37828
rect 5068 37154 5124 37156
rect 5068 37102 5070 37154
rect 5070 37102 5122 37154
rect 5122 37102 5124 37154
rect 5068 37100 5124 37102
rect 4620 36988 4676 37044
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 1820 35868 1876 35924
rect 4844 35922 4900 35924
rect 4844 35870 4846 35922
rect 4846 35870 4898 35922
rect 4898 35870 4900 35922
rect 4844 35868 4900 35870
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 5068 35084 5124 35140
rect 2492 34802 2548 34804
rect 2492 34750 2494 34802
rect 2494 34750 2546 34802
rect 2546 34750 2548 34802
rect 2492 34748 2548 34750
rect 5068 34524 5124 34580
rect 5852 38108 5908 38164
rect 6076 38050 6132 38052
rect 6076 37998 6078 38050
rect 6078 37998 6130 38050
rect 6130 37998 6132 38050
rect 6076 37996 6132 37998
rect 5964 37938 6020 37940
rect 5964 37886 5966 37938
rect 5966 37886 6018 37938
rect 6018 37886 6020 37938
rect 5964 37884 6020 37886
rect 6524 39506 6580 39508
rect 6524 39454 6526 39506
rect 6526 39454 6578 39506
rect 6578 39454 6580 39506
rect 6524 39452 6580 39454
rect 8428 39842 8484 39844
rect 8428 39790 8430 39842
rect 8430 39790 8482 39842
rect 8482 39790 8484 39842
rect 8428 39788 8484 39790
rect 9548 39788 9604 39844
rect 8092 39506 8148 39508
rect 8092 39454 8094 39506
rect 8094 39454 8146 39506
rect 8146 39454 8148 39506
rect 8092 39452 8148 39454
rect 7196 39340 7252 39396
rect 6300 39228 6356 39284
rect 7980 39004 8036 39060
rect 8316 39394 8372 39396
rect 8316 39342 8318 39394
rect 8318 39342 8370 39394
rect 8370 39342 8372 39394
rect 8316 39340 8372 39342
rect 8316 39004 8372 39060
rect 6300 38220 6356 38276
rect 6412 38556 6468 38612
rect 6076 37772 6132 37828
rect 5516 37436 5572 37492
rect 6412 37436 6468 37492
rect 6076 37266 6132 37268
rect 6076 37214 6078 37266
rect 6078 37214 6130 37266
rect 6130 37214 6132 37266
rect 6076 37212 6132 37214
rect 5964 36652 6020 36708
rect 6076 36316 6132 36372
rect 5404 35084 5460 35140
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4620 32844 4676 32900
rect 2492 32450 2548 32452
rect 2492 32398 2494 32450
rect 2494 32398 2546 32450
rect 2546 32398 2548 32450
rect 2492 32396 2548 32398
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 1708 31836 1764 31892
rect 4844 31890 4900 31892
rect 4844 31838 4846 31890
rect 4846 31838 4898 31890
rect 4898 31838 4900 31890
rect 4844 31836 4900 31838
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4956 29986 5012 29988
rect 4956 29934 4958 29986
rect 4958 29934 5010 29986
rect 5010 29934 5012 29986
rect 4956 29932 5012 29934
rect 2828 29260 2884 29316
rect 4620 29148 4676 29204
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 2604 28588 2660 28644
rect 3276 28642 3332 28644
rect 3276 28590 3278 28642
rect 3278 28590 3330 28642
rect 3330 28590 3332 28642
rect 3276 28588 3332 28590
rect 4732 28812 4788 28868
rect 5180 34076 5236 34132
rect 5740 34802 5796 34804
rect 5740 34750 5742 34802
rect 5742 34750 5794 34802
rect 5794 34750 5796 34802
rect 5740 34748 5796 34750
rect 7196 37884 7252 37940
rect 6524 37100 6580 37156
rect 5740 33346 5796 33348
rect 5740 33294 5742 33346
rect 5742 33294 5794 33346
rect 5794 33294 5796 33346
rect 5740 33292 5796 33294
rect 5292 32674 5348 32676
rect 5292 32622 5294 32674
rect 5294 32622 5346 32674
rect 5346 32622 5348 32674
rect 5292 32620 5348 32622
rect 5404 32450 5460 32452
rect 5404 32398 5406 32450
rect 5406 32398 5458 32450
rect 5458 32398 5460 32450
rect 5404 32396 5460 32398
rect 5964 33068 6020 33124
rect 6972 36988 7028 37044
rect 6972 34860 7028 34916
rect 7420 37436 7476 37492
rect 7868 37548 7924 37604
rect 9324 39618 9380 39620
rect 9324 39566 9326 39618
rect 9326 39566 9378 39618
rect 9378 39566 9380 39618
rect 9324 39564 9380 39566
rect 9772 39676 9828 39732
rect 9436 39506 9492 39508
rect 9436 39454 9438 39506
rect 9438 39454 9490 39506
rect 9490 39454 9492 39506
rect 9436 39452 9492 39454
rect 9884 39228 9940 39284
rect 10220 39564 10276 39620
rect 9772 39004 9828 39060
rect 10668 39506 10724 39508
rect 10668 39454 10670 39506
rect 10670 39454 10722 39506
rect 10722 39454 10724 39506
rect 10668 39452 10724 39454
rect 9772 38834 9828 38836
rect 9772 38782 9774 38834
rect 9774 38782 9826 38834
rect 9826 38782 9828 38834
rect 9772 38780 9828 38782
rect 8988 38556 9044 38612
rect 8316 37100 8372 37156
rect 8316 36428 8372 36484
rect 8540 35196 8596 35252
rect 7196 34300 7252 34356
rect 8092 34300 8148 34356
rect 6412 33292 6468 33348
rect 6412 32844 6468 32900
rect 6636 33122 6692 33124
rect 6636 33070 6638 33122
rect 6638 33070 6690 33122
rect 6690 33070 6692 33122
rect 6636 33068 6692 33070
rect 5852 32562 5908 32564
rect 5852 32510 5854 32562
rect 5854 32510 5906 32562
rect 5906 32510 5908 32562
rect 5852 32508 5908 32510
rect 6076 32674 6132 32676
rect 6076 32622 6078 32674
rect 6078 32622 6130 32674
rect 6130 32622 6132 32674
rect 6076 32620 6132 32622
rect 5964 31612 6020 31668
rect 5628 31500 5684 31556
rect 5292 29596 5348 29652
rect 6188 31500 6244 31556
rect 6300 31388 6356 31444
rect 6748 32732 6804 32788
rect 7084 32508 7140 32564
rect 7980 32508 8036 32564
rect 8316 32956 8372 33012
rect 8316 32732 8372 32788
rect 6524 31724 6580 31780
rect 5628 30828 5684 30884
rect 5292 29314 5348 29316
rect 5292 29262 5294 29314
rect 5294 29262 5346 29314
rect 5346 29262 5348 29314
rect 5292 29260 5348 29262
rect 6412 30882 6468 30884
rect 6412 30830 6414 30882
rect 6414 30830 6466 30882
rect 6466 30830 6468 30882
rect 6412 30828 6468 30830
rect 6076 29538 6132 29540
rect 6076 29486 6078 29538
rect 6078 29486 6130 29538
rect 6130 29486 6132 29538
rect 6076 29484 6132 29486
rect 5740 28866 5796 28868
rect 5740 28814 5742 28866
rect 5742 28814 5794 28866
rect 5794 28814 5796 28866
rect 5740 28812 5796 28814
rect 2492 26460 2548 26516
rect 1820 23548 1876 23604
rect 4956 27804 5012 27860
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 5628 27970 5684 27972
rect 5628 27918 5630 27970
rect 5630 27918 5682 27970
rect 5682 27918 5684 27970
rect 5628 27916 5684 27918
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 4396 25340 4452 25396
rect 2828 23660 2884 23716
rect 4732 24834 4788 24836
rect 4732 24782 4734 24834
rect 4734 24782 4786 24834
rect 4786 24782 4788 24834
rect 4732 24780 4788 24782
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4508 24108 4564 24164
rect 5404 26178 5460 26180
rect 5404 26126 5406 26178
rect 5406 26126 5458 26178
rect 5458 26126 5460 26178
rect 5404 26124 5460 26126
rect 6188 28364 6244 28420
rect 6188 27298 6244 27300
rect 6188 27246 6190 27298
rect 6190 27246 6242 27298
rect 6242 27246 6244 27298
rect 6188 27244 6244 27246
rect 6412 27804 6468 27860
rect 5964 26460 6020 26516
rect 7532 31724 7588 31780
rect 6748 31666 6804 31668
rect 6748 31614 6750 31666
rect 6750 31614 6802 31666
rect 6802 31614 6804 31666
rect 6748 31612 6804 31614
rect 6860 31388 6916 31444
rect 6972 30994 7028 30996
rect 6972 30942 6974 30994
rect 6974 30942 7026 30994
rect 7026 30942 7028 30994
rect 6972 30940 7028 30942
rect 7084 30716 7140 30772
rect 6860 29148 6916 29204
rect 6748 27244 6804 27300
rect 7308 29650 7364 29652
rect 7308 29598 7310 29650
rect 7310 29598 7362 29650
rect 7362 29598 7364 29650
rect 7308 29596 7364 29598
rect 8092 30940 8148 30996
rect 7308 29260 7364 29316
rect 7420 27858 7476 27860
rect 7420 27806 7422 27858
rect 7422 27806 7474 27858
rect 7474 27806 7476 27858
rect 7420 27804 7476 27806
rect 5404 24834 5460 24836
rect 5404 24782 5406 24834
rect 5406 24782 5458 24834
rect 5458 24782 5460 24834
rect 5404 24780 5460 24782
rect 5180 24556 5236 24612
rect 6412 25282 6468 25284
rect 6412 25230 6414 25282
rect 6414 25230 6466 25282
rect 6466 25230 6468 25282
rect 6412 25228 6468 25230
rect 6076 24220 6132 24276
rect 5068 23548 5124 23604
rect 5516 23548 5572 23604
rect 4956 23436 5012 23492
rect 5404 23378 5460 23380
rect 5404 23326 5406 23378
rect 5406 23326 5458 23378
rect 5458 23326 5460 23378
rect 5404 23324 5460 23326
rect 4956 23266 5012 23268
rect 4956 23214 4958 23266
rect 4958 23214 5010 23266
rect 5010 23214 5012 23266
rect 4956 23212 5012 23214
rect 5068 22930 5124 22932
rect 5068 22878 5070 22930
rect 5070 22878 5122 22930
rect 5122 22878 5124 22930
rect 5068 22876 5124 22878
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 2492 22092 2548 22148
rect 4620 21756 4676 21812
rect 5292 21810 5348 21812
rect 5292 21758 5294 21810
rect 5294 21758 5346 21810
rect 5346 21758 5348 21810
rect 5292 21756 5348 21758
rect 8204 29484 8260 29540
rect 8540 32396 8596 32452
rect 8204 27916 8260 27972
rect 6076 23772 6132 23828
rect 5964 23714 6020 23716
rect 5964 23662 5966 23714
rect 5966 23662 6018 23714
rect 6018 23662 6020 23714
rect 5964 23660 6020 23662
rect 5852 23436 5908 23492
rect 6524 23436 6580 23492
rect 6188 23266 6244 23268
rect 6188 23214 6190 23266
rect 6190 23214 6242 23266
rect 6242 23214 6244 23266
rect 6188 23212 6244 23214
rect 6412 23212 6468 23268
rect 5628 22876 5684 22932
rect 5964 22204 6020 22260
rect 6636 22258 6692 22260
rect 6636 22206 6638 22258
rect 6638 22206 6690 22258
rect 6690 22206 6692 22258
rect 6636 22204 6692 22206
rect 7756 26460 7812 26516
rect 7756 25676 7812 25732
rect 7980 25676 8036 25732
rect 7196 25394 7252 25396
rect 7196 25342 7198 25394
rect 7198 25342 7250 25394
rect 7250 25342 7252 25394
rect 7196 25340 7252 25342
rect 5740 22146 5796 22148
rect 5740 22094 5742 22146
rect 5742 22094 5794 22146
rect 5794 22094 5796 22146
rect 5740 22092 5796 22094
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 7308 25228 7364 25284
rect 7196 23436 7252 23492
rect 8204 25394 8260 25396
rect 8204 25342 8206 25394
rect 8206 25342 8258 25394
rect 8258 25342 8260 25394
rect 8204 25340 8260 25342
rect 7644 24780 7700 24836
rect 8204 23884 8260 23940
rect 8428 26290 8484 26292
rect 8428 26238 8430 26290
rect 8430 26238 8482 26290
rect 8482 26238 8484 26290
rect 8428 26236 8484 26238
rect 8876 37660 8932 37716
rect 8764 37266 8820 37268
rect 8764 37214 8766 37266
rect 8766 37214 8818 37266
rect 8818 37214 8820 37266
rect 8764 37212 8820 37214
rect 9324 37212 9380 37268
rect 9100 36370 9156 36372
rect 9100 36318 9102 36370
rect 9102 36318 9154 36370
rect 9154 36318 9156 36370
rect 9100 36316 9156 36318
rect 8876 34300 8932 34356
rect 8764 32956 8820 33012
rect 8876 32844 8932 32900
rect 8652 31612 8708 31668
rect 8652 30380 8708 30436
rect 8876 30940 8932 30996
rect 9884 37826 9940 37828
rect 9884 37774 9886 37826
rect 9886 37774 9938 37826
rect 9938 37774 9940 37826
rect 9884 37772 9940 37774
rect 10444 37772 10500 37828
rect 9548 37660 9604 37716
rect 11788 43650 11844 43652
rect 11788 43598 11790 43650
rect 11790 43598 11842 43650
rect 11842 43598 11844 43650
rect 11788 43596 11844 43598
rect 11452 43484 11508 43540
rect 13132 46674 13188 46676
rect 13132 46622 13134 46674
rect 13134 46622 13186 46674
rect 13186 46622 13188 46674
rect 13132 46620 13188 46622
rect 12796 46562 12852 46564
rect 12796 46510 12798 46562
rect 12798 46510 12850 46562
rect 12850 46510 12852 46562
rect 12796 46508 12852 46510
rect 13132 45948 13188 46004
rect 13356 46508 13412 46564
rect 12460 45666 12516 45668
rect 12460 45614 12462 45666
rect 12462 45614 12514 45666
rect 12514 45614 12516 45666
rect 12460 45612 12516 45614
rect 12236 45388 12292 45444
rect 12348 45500 12404 45556
rect 12124 45164 12180 45220
rect 13580 45388 13636 45444
rect 14028 45890 14084 45892
rect 14028 45838 14030 45890
rect 14030 45838 14082 45890
rect 14082 45838 14084 45890
rect 14028 45836 14084 45838
rect 13916 45500 13972 45556
rect 14252 46002 14308 46004
rect 14252 45950 14254 46002
rect 14254 45950 14306 46002
rect 14306 45950 14308 46002
rect 14252 45948 14308 45950
rect 14588 45836 14644 45892
rect 14252 45612 14308 45668
rect 14140 45052 14196 45108
rect 12012 43426 12068 43428
rect 12012 43374 12014 43426
rect 12014 43374 12066 43426
rect 12066 43374 12068 43426
rect 12012 43372 12068 43374
rect 12236 42866 12292 42868
rect 12236 42814 12238 42866
rect 12238 42814 12290 42866
rect 12290 42814 12292 42866
rect 12236 42812 12292 42814
rect 12684 43260 12740 43316
rect 12572 42588 12628 42644
rect 12460 40236 12516 40292
rect 12796 39730 12852 39732
rect 12796 39678 12798 39730
rect 12798 39678 12850 39730
rect 12850 39678 12852 39730
rect 12796 39676 12852 39678
rect 10780 37548 10836 37604
rect 11004 39228 11060 39284
rect 10220 37266 10276 37268
rect 10220 37214 10222 37266
rect 10222 37214 10274 37266
rect 10274 37214 10276 37266
rect 10220 37212 10276 37214
rect 9660 36988 9716 37044
rect 9436 36482 9492 36484
rect 9436 36430 9438 36482
rect 9438 36430 9490 36482
rect 9490 36430 9492 36482
rect 9436 36428 9492 36430
rect 11788 37266 11844 37268
rect 11788 37214 11790 37266
rect 11790 37214 11842 37266
rect 11842 37214 11844 37266
rect 11788 37212 11844 37214
rect 11004 37100 11060 37156
rect 10892 35868 10948 35924
rect 14028 43650 14084 43652
rect 14028 43598 14030 43650
rect 14030 43598 14082 43650
rect 14082 43598 14084 43650
rect 14028 43596 14084 43598
rect 15932 45612 15988 45668
rect 15148 45500 15204 45556
rect 16380 45500 16436 45556
rect 18060 49810 18116 49812
rect 18060 49758 18062 49810
rect 18062 49758 18114 49810
rect 18114 49758 18116 49810
rect 18060 49756 18116 49758
rect 18396 48914 18452 48916
rect 18396 48862 18398 48914
rect 18398 48862 18450 48914
rect 18450 48862 18452 48914
rect 18396 48860 18452 48862
rect 18508 48412 18564 48468
rect 17388 47404 17444 47460
rect 19836 50202 19892 50204
rect 19836 50150 19838 50202
rect 19838 50150 19890 50202
rect 19890 50150 19892 50202
rect 19836 50148 19892 50150
rect 19940 50202 19996 50204
rect 19940 50150 19942 50202
rect 19942 50150 19994 50202
rect 19994 50150 19996 50202
rect 19940 50148 19996 50150
rect 20044 50202 20100 50204
rect 20044 50150 20046 50202
rect 20046 50150 20098 50202
rect 20098 50150 20100 50202
rect 20044 50148 20100 50150
rect 22764 50316 22820 50372
rect 18956 49644 19012 49700
rect 19292 49756 19348 49812
rect 19628 49698 19684 49700
rect 19628 49646 19630 49698
rect 19630 49646 19682 49698
rect 19682 49646 19684 49698
rect 19628 49644 19684 49646
rect 20076 49644 20132 49700
rect 19628 49026 19684 49028
rect 19628 48974 19630 49026
rect 19630 48974 19682 49026
rect 19682 48974 19684 49026
rect 19628 48972 19684 48974
rect 19516 48860 19572 48916
rect 19404 48802 19460 48804
rect 19404 48750 19406 48802
rect 19406 48750 19458 48802
rect 19458 48750 19460 48802
rect 19404 48748 19460 48750
rect 20300 48914 20356 48916
rect 20300 48862 20302 48914
rect 20302 48862 20354 48914
rect 20354 48862 20356 48914
rect 20300 48860 20356 48862
rect 20188 48802 20244 48804
rect 20188 48750 20190 48802
rect 20190 48750 20242 48802
rect 20242 48750 20244 48802
rect 20188 48748 20244 48750
rect 19836 48634 19892 48636
rect 19836 48582 19838 48634
rect 19838 48582 19890 48634
rect 19890 48582 19892 48634
rect 19836 48580 19892 48582
rect 19940 48634 19996 48636
rect 19940 48582 19942 48634
rect 19942 48582 19994 48634
rect 19994 48582 19996 48634
rect 19940 48580 19996 48582
rect 20044 48634 20100 48636
rect 20044 48582 20046 48634
rect 20046 48582 20098 48634
rect 20098 48582 20100 48634
rect 20044 48580 20100 48582
rect 19404 48188 19460 48244
rect 19292 47964 19348 48020
rect 18732 46172 18788 46228
rect 16492 45612 16548 45668
rect 16268 45388 16324 45444
rect 15372 44994 15428 44996
rect 15372 44942 15374 44994
rect 15374 44942 15426 44994
rect 15426 44942 15428 44994
rect 15372 44940 15428 44942
rect 14476 44156 14532 44212
rect 14028 43036 14084 43092
rect 13020 42812 13076 42868
rect 13804 42642 13860 42644
rect 13804 42590 13806 42642
rect 13806 42590 13858 42642
rect 13858 42590 13860 42642
rect 13804 42588 13860 42590
rect 14476 42588 14532 42644
rect 14140 42194 14196 42196
rect 14140 42142 14142 42194
rect 14142 42142 14194 42194
rect 14194 42142 14196 42194
rect 14140 42140 14196 42142
rect 14588 43036 14644 43092
rect 14812 43036 14868 43092
rect 16156 44322 16212 44324
rect 16156 44270 16158 44322
rect 16158 44270 16210 44322
rect 16210 44270 16212 44322
rect 16156 44268 16212 44270
rect 14924 42642 14980 42644
rect 14924 42590 14926 42642
rect 14926 42590 14978 42642
rect 14978 42590 14980 42642
rect 14924 42588 14980 42590
rect 15148 42530 15204 42532
rect 15148 42478 15150 42530
rect 15150 42478 15202 42530
rect 15202 42478 15204 42530
rect 15148 42476 15204 42478
rect 14588 42082 14644 42084
rect 14588 42030 14590 42082
rect 14590 42030 14642 42082
rect 14642 42030 14644 42082
rect 14588 42028 14644 42030
rect 14812 42252 14868 42308
rect 15036 42194 15092 42196
rect 15036 42142 15038 42194
rect 15038 42142 15090 42194
rect 15090 42142 15092 42194
rect 15036 42140 15092 42142
rect 15148 42082 15204 42084
rect 15148 42030 15150 42082
rect 15150 42030 15202 42082
rect 15202 42030 15204 42082
rect 15148 42028 15204 42030
rect 14700 41186 14756 41188
rect 14700 41134 14702 41186
rect 14702 41134 14754 41186
rect 14754 41134 14756 41186
rect 14700 41132 14756 41134
rect 15148 40908 15204 40964
rect 16380 41916 16436 41972
rect 15372 41132 15428 41188
rect 16604 44492 16660 44548
rect 16940 45500 16996 45556
rect 16828 44322 16884 44324
rect 16828 44270 16830 44322
rect 16830 44270 16882 44322
rect 16882 44270 16884 44322
rect 16828 44268 16884 44270
rect 15596 40962 15652 40964
rect 15596 40910 15598 40962
rect 15598 40910 15650 40962
rect 15650 40910 15652 40962
rect 15596 40908 15652 40910
rect 15260 40236 15316 40292
rect 15148 39676 15204 39732
rect 13580 39618 13636 39620
rect 13580 39566 13582 39618
rect 13582 39566 13634 39618
rect 13634 39566 13636 39618
rect 13580 39564 13636 39566
rect 13468 37100 13524 37156
rect 14364 37154 14420 37156
rect 14364 37102 14366 37154
rect 14366 37102 14418 37154
rect 14418 37102 14420 37154
rect 14364 37100 14420 37102
rect 13916 36988 13972 37044
rect 12908 36428 12964 36484
rect 15484 39676 15540 39732
rect 16716 40348 16772 40404
rect 16380 39730 16436 39732
rect 16380 39678 16382 39730
rect 16382 39678 16434 39730
rect 16434 39678 16436 39730
rect 16380 39676 16436 39678
rect 16716 39564 16772 39620
rect 20412 48354 20468 48356
rect 20412 48302 20414 48354
rect 20414 48302 20466 48354
rect 20466 48302 20468 48354
rect 20412 48300 20468 48302
rect 20636 48524 20692 48580
rect 21532 48466 21588 48468
rect 21532 48414 21534 48466
rect 21534 48414 21586 48466
rect 21586 48414 21588 48466
rect 21532 48412 21588 48414
rect 22204 48466 22260 48468
rect 22204 48414 22206 48466
rect 22206 48414 22258 48466
rect 22258 48414 22260 48466
rect 22204 48412 22260 48414
rect 19740 48018 19796 48020
rect 19740 47966 19742 48018
rect 19742 47966 19794 48018
rect 19794 47966 19796 48018
rect 19740 47964 19796 47966
rect 22092 48354 22148 48356
rect 22092 48302 22094 48354
rect 22094 48302 22146 48354
rect 22146 48302 22148 48354
rect 22092 48300 22148 48302
rect 22316 48354 22372 48356
rect 22316 48302 22318 48354
rect 22318 48302 22370 48354
rect 22370 48302 22372 48354
rect 22316 48300 22372 48302
rect 21644 48242 21700 48244
rect 21644 48190 21646 48242
rect 21646 48190 21698 48242
rect 21698 48190 21700 48242
rect 21644 48188 21700 48190
rect 22652 48242 22708 48244
rect 22652 48190 22654 48242
rect 22654 48190 22706 48242
rect 22706 48190 22708 48242
rect 22652 48188 22708 48190
rect 21420 48130 21476 48132
rect 21420 48078 21422 48130
rect 21422 48078 21474 48130
rect 21474 48078 21476 48130
rect 21420 48076 21476 48078
rect 21308 47964 21364 48020
rect 19836 47066 19892 47068
rect 19836 47014 19838 47066
rect 19838 47014 19890 47066
rect 19890 47014 19892 47066
rect 19836 47012 19892 47014
rect 19940 47066 19996 47068
rect 19940 47014 19942 47066
rect 19942 47014 19994 47066
rect 19994 47014 19996 47066
rect 19940 47012 19996 47014
rect 20044 47066 20100 47068
rect 20044 47014 20046 47066
rect 20046 47014 20098 47066
rect 20098 47014 20100 47066
rect 20044 47012 20100 47014
rect 19404 46620 19460 46676
rect 19180 45666 19236 45668
rect 19180 45614 19182 45666
rect 19182 45614 19234 45666
rect 19234 45614 19236 45666
rect 19180 45612 19236 45614
rect 18620 45276 18676 45332
rect 18060 45218 18116 45220
rect 18060 45166 18062 45218
rect 18062 45166 18114 45218
rect 18114 45166 18116 45218
rect 18060 45164 18116 45166
rect 18844 45164 18900 45220
rect 18284 45106 18340 45108
rect 18284 45054 18286 45106
rect 18286 45054 18338 45106
rect 18338 45054 18340 45106
rect 18284 45052 18340 45054
rect 19068 45218 19124 45220
rect 19068 45166 19070 45218
rect 19070 45166 19122 45218
rect 19122 45166 19124 45218
rect 19068 45164 19124 45166
rect 19068 44882 19124 44884
rect 19068 44830 19070 44882
rect 19070 44830 19122 44882
rect 19122 44830 19124 44882
rect 19068 44828 19124 44830
rect 18284 44604 18340 44660
rect 17276 44546 17332 44548
rect 17276 44494 17278 44546
rect 17278 44494 17330 44546
rect 17330 44494 17332 44546
rect 17276 44492 17332 44494
rect 17724 44434 17780 44436
rect 17724 44382 17726 44434
rect 17726 44382 17778 44434
rect 17778 44382 17780 44434
rect 17724 44380 17780 44382
rect 18172 44322 18228 44324
rect 18172 44270 18174 44322
rect 18174 44270 18226 44322
rect 18226 44270 18228 44322
rect 18172 44268 18228 44270
rect 18396 44380 18452 44436
rect 17052 43372 17108 43428
rect 18620 44434 18676 44436
rect 18620 44382 18622 44434
rect 18622 44382 18674 44434
rect 18674 44382 18676 44434
rect 18620 44380 18676 44382
rect 21084 46898 21140 46900
rect 21084 46846 21086 46898
rect 21086 46846 21138 46898
rect 21138 46846 21140 46898
rect 21084 46844 21140 46846
rect 20412 46786 20468 46788
rect 20412 46734 20414 46786
rect 20414 46734 20466 46786
rect 20466 46734 20468 46786
rect 20412 46732 20468 46734
rect 20972 46786 21028 46788
rect 20972 46734 20974 46786
rect 20974 46734 21026 46786
rect 21026 46734 21028 46786
rect 20972 46732 21028 46734
rect 20300 46674 20356 46676
rect 20300 46622 20302 46674
rect 20302 46622 20354 46674
rect 20354 46622 20356 46674
rect 20300 46620 20356 46622
rect 22540 46508 22596 46564
rect 22428 45890 22484 45892
rect 22428 45838 22430 45890
rect 22430 45838 22482 45890
rect 22482 45838 22484 45890
rect 22428 45836 22484 45838
rect 19836 45498 19892 45500
rect 19836 45446 19838 45498
rect 19838 45446 19890 45498
rect 19890 45446 19892 45498
rect 19836 45444 19892 45446
rect 19940 45498 19996 45500
rect 19940 45446 19942 45498
rect 19942 45446 19994 45498
rect 19994 45446 19996 45498
rect 19940 45444 19996 45446
rect 20044 45498 20100 45500
rect 20044 45446 20046 45498
rect 20046 45446 20098 45498
rect 20098 45446 20100 45498
rect 20044 45444 20100 45446
rect 22652 45500 22708 45556
rect 19628 45276 19684 45332
rect 21980 45388 22036 45444
rect 19740 44604 19796 44660
rect 19852 44828 19908 44884
rect 18396 44210 18452 44212
rect 18396 44158 18398 44210
rect 18398 44158 18450 44210
rect 18450 44158 18452 44210
rect 18396 44156 18452 44158
rect 21868 45052 21924 45108
rect 19516 44098 19572 44100
rect 19516 44046 19518 44098
rect 19518 44046 19570 44098
rect 19570 44046 19572 44098
rect 19516 44044 19572 44046
rect 18732 43708 18788 43764
rect 19292 43708 19348 43764
rect 20300 44098 20356 44100
rect 20300 44046 20302 44098
rect 20302 44046 20354 44098
rect 20354 44046 20356 44098
rect 20300 44044 20356 44046
rect 22540 44210 22596 44212
rect 22540 44158 22542 44210
rect 22542 44158 22594 44210
rect 22594 44158 22596 44210
rect 22540 44156 22596 44158
rect 22092 44098 22148 44100
rect 22092 44046 22094 44098
rect 22094 44046 22146 44098
rect 22146 44046 22148 44098
rect 22092 44044 22148 44046
rect 19836 43930 19892 43932
rect 19836 43878 19838 43930
rect 19838 43878 19890 43930
rect 19890 43878 19892 43930
rect 19836 43876 19892 43878
rect 19940 43930 19996 43932
rect 19940 43878 19942 43930
rect 19942 43878 19994 43930
rect 19994 43878 19996 43930
rect 19940 43876 19996 43878
rect 20044 43930 20100 43932
rect 20044 43878 20046 43930
rect 20046 43878 20098 43930
rect 20098 43878 20100 43930
rect 20044 43876 20100 43878
rect 18956 43538 19012 43540
rect 18956 43486 18958 43538
rect 18958 43486 19010 43538
rect 19010 43486 19012 43538
rect 18956 43484 19012 43486
rect 18508 43426 18564 43428
rect 18508 43374 18510 43426
rect 18510 43374 18562 43426
rect 18562 43374 18564 43426
rect 18508 43372 18564 43374
rect 18060 41356 18116 41412
rect 21420 43762 21476 43764
rect 21420 43710 21422 43762
rect 21422 43710 21474 43762
rect 21474 43710 21476 43762
rect 21420 43708 21476 43710
rect 19836 42362 19892 42364
rect 19836 42310 19838 42362
rect 19838 42310 19890 42362
rect 19890 42310 19892 42362
rect 19836 42308 19892 42310
rect 19940 42362 19996 42364
rect 19940 42310 19942 42362
rect 19942 42310 19994 42362
rect 19994 42310 19996 42362
rect 19940 42308 19996 42310
rect 20044 42362 20100 42364
rect 20044 42310 20046 42362
rect 20046 42310 20098 42362
rect 20098 42310 20100 42362
rect 20044 42308 20100 42310
rect 18620 40402 18676 40404
rect 18620 40350 18622 40402
rect 18622 40350 18674 40402
rect 18674 40350 18676 40402
rect 18620 40348 18676 40350
rect 19068 40402 19124 40404
rect 19068 40350 19070 40402
rect 19070 40350 19122 40402
rect 19122 40350 19124 40402
rect 19068 40348 19124 40350
rect 16604 38834 16660 38836
rect 16604 38782 16606 38834
rect 16606 38782 16658 38834
rect 16658 38782 16660 38834
rect 16604 38780 16660 38782
rect 15932 37996 15988 38052
rect 15484 36316 15540 36372
rect 11676 35868 11732 35924
rect 9548 34860 9604 34916
rect 9436 33122 9492 33124
rect 9436 33070 9438 33122
rect 9438 33070 9490 33122
rect 9490 33070 9492 33122
rect 9436 33068 9492 33070
rect 9884 33180 9940 33236
rect 9100 31778 9156 31780
rect 9100 31726 9102 31778
rect 9102 31726 9154 31778
rect 9154 31726 9156 31778
rect 9100 31724 9156 31726
rect 10556 34130 10612 34132
rect 10556 34078 10558 34130
rect 10558 34078 10610 34130
rect 10610 34078 10612 34130
rect 10556 34076 10612 34078
rect 11116 34076 11172 34132
rect 14364 34914 14420 34916
rect 14364 34862 14366 34914
rect 14366 34862 14418 34914
rect 14418 34862 14420 34914
rect 14364 34860 14420 34862
rect 14812 34914 14868 34916
rect 14812 34862 14814 34914
rect 14814 34862 14866 34914
rect 14866 34862 14868 34914
rect 14812 34860 14868 34862
rect 13804 34130 13860 34132
rect 13804 34078 13806 34130
rect 13806 34078 13858 34130
rect 13858 34078 13860 34130
rect 13804 34076 13860 34078
rect 9324 31500 9380 31556
rect 9212 31052 9268 31108
rect 9884 31554 9940 31556
rect 9884 31502 9886 31554
rect 9886 31502 9938 31554
rect 9938 31502 9940 31554
rect 9884 31500 9940 31502
rect 10668 33234 10724 33236
rect 10668 33182 10670 33234
rect 10670 33182 10722 33234
rect 10722 33182 10724 33234
rect 10668 33180 10724 33182
rect 10220 33122 10276 33124
rect 10220 33070 10222 33122
rect 10222 33070 10274 33122
rect 10274 33070 10276 33122
rect 10220 33068 10276 33070
rect 13020 32450 13076 32452
rect 13020 32398 13022 32450
rect 13022 32398 13074 32450
rect 13074 32398 13076 32450
rect 13020 32396 13076 32398
rect 10556 31948 10612 32004
rect 13692 32396 13748 32452
rect 13356 31948 13412 32004
rect 11116 31890 11172 31892
rect 11116 31838 11118 31890
rect 11118 31838 11170 31890
rect 11170 31838 11172 31890
rect 11116 31836 11172 31838
rect 10108 31052 10164 31108
rect 9548 30434 9604 30436
rect 9548 30382 9550 30434
rect 9550 30382 9602 30434
rect 9602 30382 9604 30434
rect 9548 30380 9604 30382
rect 9772 30322 9828 30324
rect 9772 30270 9774 30322
rect 9774 30270 9826 30322
rect 9826 30270 9828 30322
rect 9772 30268 9828 30270
rect 10220 30268 10276 30324
rect 10108 29932 10164 29988
rect 10556 31106 10612 31108
rect 10556 31054 10558 31106
rect 10558 31054 10610 31106
rect 10610 31054 10612 31106
rect 10556 31052 10612 31054
rect 10668 30268 10724 30324
rect 8988 28364 9044 28420
rect 8988 27020 9044 27076
rect 8540 25676 8596 25732
rect 8876 26908 8932 26964
rect 8428 25228 8484 25284
rect 9772 27020 9828 27076
rect 14364 32562 14420 32564
rect 14364 32510 14366 32562
rect 14366 32510 14418 32562
rect 14418 32510 14420 32562
rect 14364 32508 14420 32510
rect 14588 31890 14644 31892
rect 14588 31838 14590 31890
rect 14590 31838 14642 31890
rect 14642 31838 14644 31890
rect 14588 31836 14644 31838
rect 13580 31500 13636 31556
rect 13356 30156 13412 30212
rect 13468 30268 13524 30324
rect 14140 30940 14196 30996
rect 11340 28588 11396 28644
rect 11900 28642 11956 28644
rect 11900 28590 11902 28642
rect 11902 28590 11954 28642
rect 11954 28590 11956 28642
rect 11900 28588 11956 28590
rect 11564 28082 11620 28084
rect 11564 28030 11566 28082
rect 11566 28030 11618 28082
rect 11618 28030 11620 28082
rect 11564 28028 11620 28030
rect 12684 28028 12740 28084
rect 9996 26962 10052 26964
rect 9996 26910 9998 26962
rect 9998 26910 10050 26962
rect 10050 26910 10052 26962
rect 9996 26908 10052 26910
rect 9548 26236 9604 26292
rect 8652 25340 8708 25396
rect 7644 23266 7700 23268
rect 7644 23214 7646 23266
rect 7646 23214 7698 23266
rect 7698 23214 7700 23266
rect 7644 23212 7700 23214
rect 8316 23714 8372 23716
rect 8316 23662 8318 23714
rect 8318 23662 8370 23714
rect 8370 23662 8372 23714
rect 8316 23660 8372 23662
rect 8540 23884 8596 23940
rect 7420 23042 7476 23044
rect 7420 22990 7422 23042
rect 7422 22990 7474 23042
rect 7474 22990 7476 23042
rect 7420 22988 7476 22990
rect 8092 21810 8148 21812
rect 8092 21758 8094 21810
rect 8094 21758 8146 21810
rect 8146 21758 8148 21810
rect 8092 21756 8148 21758
rect 8876 23938 8932 23940
rect 8876 23886 8878 23938
rect 8878 23886 8930 23938
rect 8930 23886 8932 23938
rect 8876 23884 8932 23886
rect 8764 23826 8820 23828
rect 8764 23774 8766 23826
rect 8766 23774 8818 23826
rect 8818 23774 8820 23826
rect 8764 23772 8820 23774
rect 9660 25452 9716 25508
rect 11004 27970 11060 27972
rect 11004 27918 11006 27970
rect 11006 27918 11058 27970
rect 11058 27918 11060 27970
rect 11004 27916 11060 27918
rect 11564 27132 11620 27188
rect 11116 27074 11172 27076
rect 11116 27022 11118 27074
rect 11118 27022 11170 27074
rect 11170 27022 11172 27074
rect 11116 27020 11172 27022
rect 10780 26908 10836 26964
rect 14812 32562 14868 32564
rect 14812 32510 14814 32562
rect 14814 32510 14866 32562
rect 14866 32510 14868 32562
rect 14812 32508 14868 32510
rect 15484 34690 15540 34692
rect 15484 34638 15486 34690
rect 15486 34638 15538 34690
rect 15538 34638 15540 34690
rect 15484 34636 15540 34638
rect 15036 33346 15092 33348
rect 15036 33294 15038 33346
rect 15038 33294 15090 33346
rect 15090 33294 15092 33346
rect 15036 33292 15092 33294
rect 15036 32956 15092 33012
rect 16268 36988 16324 37044
rect 16044 36370 16100 36372
rect 16044 36318 16046 36370
rect 16046 36318 16098 36370
rect 16098 36318 16100 36370
rect 16044 36316 16100 36318
rect 15484 33516 15540 33572
rect 15372 32956 15428 33012
rect 16156 32674 16212 32676
rect 16156 32622 16158 32674
rect 16158 32622 16210 32674
rect 16210 32622 16212 32674
rect 16156 32620 16212 32622
rect 16604 35586 16660 35588
rect 16604 35534 16606 35586
rect 16606 35534 16658 35586
rect 16658 35534 16660 35586
rect 16604 35532 16660 35534
rect 16604 34636 16660 34692
rect 16828 38332 16884 38388
rect 19516 41580 19572 41636
rect 16604 32732 16660 32788
rect 14812 29596 14868 29652
rect 11788 27186 11844 27188
rect 11788 27134 11790 27186
rect 11790 27134 11842 27186
rect 11842 27134 11844 27186
rect 11788 27132 11844 27134
rect 14700 27020 14756 27076
rect 11676 26908 11732 26964
rect 9100 23714 9156 23716
rect 9100 23662 9102 23714
rect 9102 23662 9154 23714
rect 9154 23662 9156 23714
rect 9100 23660 9156 23662
rect 8428 22988 8484 23044
rect 8988 23042 9044 23044
rect 8988 22990 8990 23042
rect 8990 22990 9042 23042
rect 9042 22990 9044 23042
rect 8988 22988 9044 22990
rect 8876 22930 8932 22932
rect 8876 22878 8878 22930
rect 8878 22878 8930 22930
rect 8930 22878 8932 22930
rect 8876 22876 8932 22878
rect 8652 21756 8708 21812
rect 7084 20076 7140 20132
rect 4956 19852 5012 19908
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 6412 19852 6468 19908
rect 8652 20412 8708 20468
rect 8764 20636 8820 20692
rect 7084 19740 7140 19796
rect 4956 19010 5012 19012
rect 4956 18958 4958 19010
rect 4958 18958 5010 19010
rect 5010 18958 5012 19010
rect 4956 18956 5012 18958
rect 2492 18450 2548 18452
rect 2492 18398 2494 18450
rect 2494 18398 2546 18450
rect 2546 18398 2548 18450
rect 2492 18396 2548 18398
rect 4620 18338 4676 18340
rect 4620 18286 4622 18338
rect 4622 18286 4674 18338
rect 4674 18286 4676 18338
rect 4620 18284 4676 18286
rect 5628 18956 5684 19012
rect 6188 19010 6244 19012
rect 6188 18958 6190 19010
rect 6190 18958 6242 19010
rect 6242 18958 6244 19010
rect 6188 18956 6244 18958
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 5516 18284 5572 18340
rect 5516 17500 5572 17556
rect 1820 16828 1876 16884
rect 5068 16828 5124 16884
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 2604 15314 2660 15316
rect 2604 15262 2606 15314
rect 2606 15262 2658 15314
rect 2658 15262 2660 15314
rect 2604 15260 2660 15262
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 6412 17724 6468 17780
rect 6636 18844 6692 18900
rect 7644 19740 7700 19796
rect 7084 19068 7140 19124
rect 6300 17554 6356 17556
rect 6300 17502 6302 17554
rect 6302 17502 6354 17554
rect 6354 17502 6356 17554
rect 6300 17500 6356 17502
rect 6188 16098 6244 16100
rect 6188 16046 6190 16098
rect 6190 16046 6242 16098
rect 6242 16046 6244 16098
rect 6188 16044 6244 16046
rect 4956 15426 5012 15428
rect 4956 15374 4958 15426
rect 4958 15374 5010 15426
rect 5010 15374 5012 15426
rect 4956 15372 5012 15374
rect 2492 13580 2548 13636
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4844 13244 4900 13300
rect 6188 14252 6244 14308
rect 4956 13074 5012 13076
rect 4956 13022 4958 13074
rect 4958 13022 5010 13074
rect 5010 13022 5012 13074
rect 4956 13020 5012 13022
rect 5068 12962 5124 12964
rect 5068 12910 5070 12962
rect 5070 12910 5122 12962
rect 5122 12910 5124 12962
rect 5068 12908 5124 12910
rect 4956 12796 5012 12852
rect 5740 13020 5796 13076
rect 6076 13634 6132 13636
rect 6076 13582 6078 13634
rect 6078 13582 6130 13634
rect 6130 13582 6132 13634
rect 6076 13580 6132 13582
rect 6412 16492 6468 16548
rect 7980 19292 8036 19348
rect 8652 20130 8708 20132
rect 8652 20078 8654 20130
rect 8654 20078 8706 20130
rect 8706 20078 8708 20130
rect 8652 20076 8708 20078
rect 8316 20018 8372 20020
rect 8316 19966 8318 20018
rect 8318 19966 8370 20018
rect 8370 19966 8372 20018
rect 8316 19964 8372 19966
rect 8540 19346 8596 19348
rect 8540 19294 8542 19346
rect 8542 19294 8594 19346
rect 8594 19294 8596 19346
rect 8540 19292 8596 19294
rect 8316 19068 8372 19124
rect 6972 17724 7028 17780
rect 6524 16156 6580 16212
rect 7980 17724 8036 17780
rect 7084 16044 7140 16100
rect 7084 15426 7140 15428
rect 7084 15374 7086 15426
rect 7086 15374 7138 15426
rect 7138 15374 7140 15426
rect 7084 15372 7140 15374
rect 7532 16156 7588 16212
rect 7308 16098 7364 16100
rect 7308 16046 7310 16098
rect 7310 16046 7362 16098
rect 7362 16046 7364 16098
rect 7308 16044 7364 16046
rect 9772 25004 9828 25060
rect 10668 24668 10724 24724
rect 9212 22876 9268 22932
rect 9660 21810 9716 21812
rect 9660 21758 9662 21810
rect 9662 21758 9714 21810
rect 9714 21758 9716 21810
rect 9660 21756 9716 21758
rect 10108 24610 10164 24612
rect 10108 24558 10110 24610
rect 10110 24558 10162 24610
rect 10162 24558 10164 24610
rect 10108 24556 10164 24558
rect 11116 25506 11172 25508
rect 11116 25454 11118 25506
rect 11118 25454 11170 25506
rect 11170 25454 11172 25506
rect 11116 25452 11172 25454
rect 11004 25228 11060 25284
rect 10556 23772 10612 23828
rect 9996 21868 10052 21924
rect 9996 21474 10052 21476
rect 9996 21422 9998 21474
rect 9998 21422 10050 21474
rect 10050 21422 10052 21474
rect 9996 21420 10052 21422
rect 9884 20972 9940 21028
rect 9660 20412 9716 20468
rect 8876 19740 8932 19796
rect 8988 20018 9044 20020
rect 8988 19966 8990 20018
rect 8990 19966 9042 20018
rect 9042 19966 9044 20018
rect 8988 19964 9044 19966
rect 8988 19404 9044 19460
rect 9100 19292 9156 19348
rect 8316 15372 8372 15428
rect 7532 15314 7588 15316
rect 7532 15262 7534 15314
rect 7534 15262 7586 15314
rect 7586 15262 7588 15314
rect 7532 15260 7588 15262
rect 8092 15314 8148 15316
rect 8092 15262 8094 15314
rect 8094 15262 8146 15314
rect 8146 15262 8148 15314
rect 8092 15260 8148 15262
rect 7084 14306 7140 14308
rect 7084 14254 7086 14306
rect 7086 14254 7138 14306
rect 7138 14254 7140 14306
rect 7084 14252 7140 14254
rect 6412 13916 6468 13972
rect 6412 13244 6468 13300
rect 7196 13468 7252 13524
rect 7308 13970 7364 13972
rect 7308 13918 7310 13970
rect 7310 13918 7362 13970
rect 7362 13918 7364 13970
rect 7308 13916 7364 13918
rect 8092 14252 8148 14308
rect 6188 13186 6244 13188
rect 6188 13134 6190 13186
rect 6190 13134 6242 13186
rect 6242 13134 6244 13186
rect 6188 13132 6244 13134
rect 5964 12908 6020 12964
rect 6860 12962 6916 12964
rect 6860 12910 6862 12962
rect 6862 12910 6914 12962
rect 6914 12910 6916 12962
rect 6860 12908 6916 12910
rect 5628 12850 5684 12852
rect 5628 12798 5630 12850
rect 5630 12798 5682 12850
rect 5682 12798 5684 12850
rect 5628 12796 5684 12798
rect 5964 12684 6020 12740
rect 1820 12012 1876 12068
rect 4844 12066 4900 12068
rect 4844 12014 4846 12066
rect 4846 12014 4898 12066
rect 4898 12014 4900 12066
rect 4844 12012 4900 12014
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4284 11228 4340 11284
rect 2492 11116 2548 11172
rect 4172 10780 4228 10836
rect 5852 12236 5908 12292
rect 5964 11452 6020 11508
rect 4620 10780 4676 10836
rect 5740 11170 5796 11172
rect 5740 11118 5742 11170
rect 5742 11118 5794 11170
rect 5794 11118 5796 11170
rect 5740 11116 5796 11118
rect 6636 11394 6692 11396
rect 6636 11342 6638 11394
rect 6638 11342 6690 11394
rect 6690 11342 6692 11394
rect 6636 11340 6692 11342
rect 6076 11116 6132 11172
rect 7196 13074 7252 13076
rect 7196 13022 7198 13074
rect 7198 13022 7250 13074
rect 7250 13022 7252 13074
rect 7196 13020 7252 13022
rect 6972 11170 7028 11172
rect 6972 11118 6974 11170
rect 6974 11118 7026 11170
rect 7026 11118 7028 11170
rect 6972 11116 7028 11118
rect 5068 10834 5124 10836
rect 5068 10782 5070 10834
rect 5070 10782 5122 10834
rect 5122 10782 5124 10834
rect 5068 10780 5124 10782
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 7196 10108 7252 10164
rect 4172 9772 4228 9828
rect 6972 9826 7028 9828
rect 6972 9774 6974 9826
rect 6974 9774 7026 9826
rect 7026 9774 7028 9826
rect 6972 9772 7028 9774
rect 7868 11506 7924 11508
rect 7868 11454 7870 11506
rect 7870 11454 7922 11506
rect 7922 11454 7924 11506
rect 7868 11452 7924 11454
rect 7756 10780 7812 10836
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 7644 9772 7700 9828
rect 7756 9266 7812 9268
rect 7756 9214 7758 9266
rect 7758 9214 7810 9266
rect 7810 9214 7812 9266
rect 7756 9212 7812 9214
rect 7308 8092 7364 8148
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 8092 13468 8148 13524
rect 10556 20972 10612 21028
rect 9772 19906 9828 19908
rect 9772 19854 9774 19906
rect 9774 19854 9826 19906
rect 9826 19854 9828 19906
rect 9772 19852 9828 19854
rect 10108 19740 10164 19796
rect 10108 19122 10164 19124
rect 10108 19070 10110 19122
rect 10110 19070 10162 19122
rect 10162 19070 10164 19122
rect 10108 19068 10164 19070
rect 10444 19010 10500 19012
rect 10444 18958 10446 19010
rect 10446 18958 10498 19010
rect 10498 18958 10500 19010
rect 10444 18956 10500 18958
rect 11116 24892 11172 24948
rect 11564 24668 11620 24724
rect 11116 24556 11172 24612
rect 12236 26962 12292 26964
rect 12236 26910 12238 26962
rect 12238 26910 12290 26962
rect 12290 26910 12292 26962
rect 12236 26908 12292 26910
rect 16156 30828 16212 30884
rect 15596 30716 15652 30772
rect 15372 29148 15428 29204
rect 15932 29148 15988 29204
rect 15484 27916 15540 27972
rect 16156 27858 16212 27860
rect 16156 27806 16158 27858
rect 16158 27806 16210 27858
rect 16210 27806 16212 27858
rect 16156 27804 16212 27806
rect 15148 25564 15204 25620
rect 11900 25282 11956 25284
rect 11900 25230 11902 25282
rect 11902 25230 11954 25282
rect 11954 25230 11956 25282
rect 11900 25228 11956 25230
rect 11900 24892 11956 24948
rect 14476 24722 14532 24724
rect 14476 24670 14478 24722
rect 14478 24670 14530 24722
rect 14530 24670 14532 24722
rect 14476 24668 14532 24670
rect 16156 24722 16212 24724
rect 16156 24670 16158 24722
rect 16158 24670 16210 24722
rect 16210 24670 16212 24722
rect 16156 24668 16212 24670
rect 11676 24556 11732 24612
rect 12348 24556 12404 24612
rect 15708 23938 15764 23940
rect 15708 23886 15710 23938
rect 15710 23886 15762 23938
rect 15762 23886 15764 23938
rect 15708 23884 15764 23886
rect 15372 23826 15428 23828
rect 15372 23774 15374 23826
rect 15374 23774 15426 23826
rect 15426 23774 15428 23826
rect 15372 23772 15428 23774
rect 13468 23042 13524 23044
rect 13468 22990 13470 23042
rect 13470 22990 13522 23042
rect 13522 22990 13524 23042
rect 13468 22988 13524 22990
rect 12684 21756 12740 21812
rect 11340 21644 11396 21700
rect 14028 21810 14084 21812
rect 14028 21758 14030 21810
rect 14030 21758 14082 21810
rect 14082 21758 14084 21810
rect 14028 21756 14084 21758
rect 13468 21644 13524 21700
rect 11004 20748 11060 20804
rect 15036 21308 15092 21364
rect 13804 20690 13860 20692
rect 13804 20638 13806 20690
rect 13806 20638 13858 20690
rect 13858 20638 13860 20690
rect 13804 20636 13860 20638
rect 12012 19852 12068 19908
rect 11116 19740 11172 19796
rect 11004 18956 11060 19012
rect 10556 17164 10612 17220
rect 10220 16940 10276 16996
rect 9660 16882 9716 16884
rect 9660 16830 9662 16882
rect 9662 16830 9714 16882
rect 9714 16830 9716 16882
rect 9660 16828 9716 16830
rect 9884 16492 9940 16548
rect 8764 15426 8820 15428
rect 8764 15374 8766 15426
rect 8766 15374 8818 15426
rect 8818 15374 8820 15426
rect 8764 15372 8820 15374
rect 8652 15260 8708 15316
rect 9436 15148 9492 15204
rect 9548 15260 9604 15316
rect 8316 13132 8372 13188
rect 8316 11954 8372 11956
rect 8316 11902 8318 11954
rect 8318 11902 8370 11954
rect 8370 11902 8372 11954
rect 8316 11900 8372 11902
rect 8204 11452 8260 11508
rect 8652 11282 8708 11284
rect 8652 11230 8654 11282
rect 8654 11230 8706 11282
rect 8706 11230 8708 11282
rect 8652 11228 8708 11230
rect 7868 8258 7924 8260
rect 7868 8206 7870 8258
rect 7870 8206 7922 8258
rect 7922 8206 7924 8258
rect 7868 8204 7924 8206
rect 8988 8258 9044 8260
rect 8988 8206 8990 8258
rect 8990 8206 9042 8258
rect 9042 8206 9044 8258
rect 8988 8204 9044 8206
rect 8876 8146 8932 8148
rect 8876 8094 8878 8146
rect 8878 8094 8930 8146
rect 8930 8094 8932 8146
rect 8876 8092 8932 8094
rect 8092 8034 8148 8036
rect 8092 7982 8094 8034
rect 8094 7982 8146 8034
rect 8146 7982 8148 8034
rect 8092 7980 8148 7982
rect 8316 7698 8372 7700
rect 8316 7646 8318 7698
rect 8318 7646 8370 7698
rect 8370 7646 8372 7698
rect 8316 7644 8372 7646
rect 9884 15260 9940 15316
rect 9772 15148 9828 15204
rect 10444 15036 10500 15092
rect 11452 19458 11508 19460
rect 11452 19406 11454 19458
rect 11454 19406 11506 19458
rect 11506 19406 11508 19458
rect 11452 19404 11508 19406
rect 11228 19346 11284 19348
rect 11228 19294 11230 19346
rect 11230 19294 11282 19346
rect 11282 19294 11284 19346
rect 11228 19292 11284 19294
rect 12012 19346 12068 19348
rect 12012 19294 12014 19346
rect 12014 19294 12066 19346
rect 12066 19294 12068 19346
rect 12012 19292 12068 19294
rect 15260 20690 15316 20692
rect 15260 20638 15262 20690
rect 15262 20638 15314 20690
rect 15314 20638 15316 20690
rect 15260 20636 15316 20638
rect 14364 19068 14420 19124
rect 14476 20076 14532 20132
rect 11564 17052 11620 17108
rect 11676 16940 11732 16996
rect 11900 16828 11956 16884
rect 11788 16098 11844 16100
rect 11788 16046 11790 16098
rect 11790 16046 11842 16098
rect 11842 16046 11844 16098
rect 11788 16044 11844 16046
rect 12348 17052 12404 17108
rect 13468 17164 13524 17220
rect 11900 15820 11956 15876
rect 12124 16268 12180 16324
rect 11116 15036 11172 15092
rect 11340 14530 11396 14532
rect 11340 14478 11342 14530
rect 11342 14478 11394 14530
rect 11394 14478 11396 14530
rect 11340 14476 11396 14478
rect 13132 17052 13188 17108
rect 13020 16994 13076 16996
rect 13020 16942 13022 16994
rect 13022 16942 13074 16994
rect 13074 16942 13076 16994
rect 13020 16940 13076 16942
rect 13244 16882 13300 16884
rect 13244 16830 13246 16882
rect 13246 16830 13298 16882
rect 13298 16830 13300 16882
rect 13244 16828 13300 16830
rect 14924 20018 14980 20020
rect 14924 19966 14926 20018
rect 14926 19966 14978 20018
rect 14978 19966 14980 20018
rect 14924 19964 14980 19966
rect 15484 20018 15540 20020
rect 15484 19966 15486 20018
rect 15486 19966 15538 20018
rect 15538 19966 15540 20018
rect 15484 19964 15540 19966
rect 15148 19740 15204 19796
rect 16380 20690 16436 20692
rect 16380 20638 16382 20690
rect 16382 20638 16434 20690
rect 16434 20638 16436 20690
rect 16380 20636 16436 20638
rect 15820 20130 15876 20132
rect 15820 20078 15822 20130
rect 15822 20078 15874 20130
rect 15874 20078 15876 20130
rect 15820 20076 15876 20078
rect 16940 32396 16996 32452
rect 16604 31836 16660 31892
rect 16716 30882 16772 30884
rect 16716 30830 16718 30882
rect 16718 30830 16770 30882
rect 16770 30830 16772 30882
rect 16716 30828 16772 30830
rect 16828 29260 16884 29316
rect 16604 28028 16660 28084
rect 16716 27858 16772 27860
rect 16716 27806 16718 27858
rect 16718 27806 16770 27858
rect 16770 27806 16772 27858
rect 16716 27804 16772 27806
rect 16828 27746 16884 27748
rect 16828 27694 16830 27746
rect 16830 27694 16882 27746
rect 16882 27694 16884 27746
rect 16828 27692 16884 27694
rect 16828 25340 16884 25396
rect 16716 24892 16772 24948
rect 17612 38780 17668 38836
rect 18172 38892 18228 38948
rect 19068 38332 19124 38388
rect 18060 38050 18116 38052
rect 18060 37998 18062 38050
rect 18062 37998 18114 38050
rect 18114 37998 18116 38050
rect 18060 37996 18116 37998
rect 17724 37884 17780 37940
rect 18284 36540 18340 36596
rect 19068 37266 19124 37268
rect 19068 37214 19070 37266
rect 19070 37214 19122 37266
rect 19122 37214 19124 37266
rect 19068 37212 19124 37214
rect 18732 36594 18788 36596
rect 18732 36542 18734 36594
rect 18734 36542 18786 36594
rect 18786 36542 18788 36594
rect 18732 36540 18788 36542
rect 17724 36482 17780 36484
rect 17724 36430 17726 36482
rect 17726 36430 17778 36482
rect 17778 36430 17780 36482
rect 17724 36428 17780 36430
rect 17948 33964 18004 34020
rect 17724 32396 17780 32452
rect 17836 31500 17892 31556
rect 17948 30994 18004 30996
rect 17948 30942 17950 30994
rect 17950 30942 18002 30994
rect 18002 30942 18004 30994
rect 17948 30940 18004 30942
rect 18508 35196 18564 35252
rect 19180 36482 19236 36484
rect 19180 36430 19182 36482
rect 19182 36430 19234 36482
rect 19234 36430 19236 36482
rect 19180 36428 19236 36430
rect 19836 40794 19892 40796
rect 19836 40742 19838 40794
rect 19838 40742 19890 40794
rect 19890 40742 19892 40794
rect 19836 40740 19892 40742
rect 19940 40794 19996 40796
rect 19940 40742 19942 40794
rect 19942 40742 19994 40794
rect 19994 40742 19996 40794
rect 19940 40740 19996 40742
rect 20044 40794 20100 40796
rect 20044 40742 20046 40794
rect 20046 40742 20098 40794
rect 20098 40742 20100 40794
rect 20044 40740 20100 40742
rect 19740 40514 19796 40516
rect 19740 40462 19742 40514
rect 19742 40462 19794 40514
rect 19794 40462 19796 40514
rect 19740 40460 19796 40462
rect 19628 40348 19684 40404
rect 19836 39226 19892 39228
rect 19836 39174 19838 39226
rect 19838 39174 19890 39226
rect 19890 39174 19892 39226
rect 19836 39172 19892 39174
rect 19940 39226 19996 39228
rect 19940 39174 19942 39226
rect 19942 39174 19994 39226
rect 19994 39174 19996 39226
rect 19940 39172 19996 39174
rect 20044 39226 20100 39228
rect 20044 39174 20046 39226
rect 20046 39174 20098 39226
rect 20098 39174 20100 39226
rect 20044 39172 20100 39174
rect 19740 38946 19796 38948
rect 19740 38894 19742 38946
rect 19742 38894 19794 38946
rect 19794 38894 19796 38946
rect 19740 38892 19796 38894
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 20076 36316 20132 36372
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19292 35532 19348 35588
rect 18844 34636 18900 34692
rect 18732 34242 18788 34244
rect 18732 34190 18734 34242
rect 18734 34190 18786 34242
rect 18786 34190 18788 34242
rect 18732 34188 18788 34190
rect 18284 32844 18340 32900
rect 19404 34690 19460 34692
rect 19404 34638 19406 34690
rect 19406 34638 19458 34690
rect 19458 34638 19460 34690
rect 19404 34636 19460 34638
rect 20188 34636 20244 34692
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19180 34018 19236 34020
rect 19180 33966 19182 34018
rect 19182 33966 19234 34018
rect 19234 33966 19236 34018
rect 19180 33964 19236 33966
rect 18956 33516 19012 33572
rect 19628 33404 19684 33460
rect 19404 33346 19460 33348
rect 19404 33294 19406 33346
rect 19406 33294 19458 33346
rect 19458 33294 19460 33346
rect 19404 33292 19460 33294
rect 18844 32844 18900 32900
rect 17500 29426 17556 29428
rect 17500 29374 17502 29426
rect 17502 29374 17554 29426
rect 17554 29374 17556 29426
rect 17500 29372 17556 29374
rect 17276 28642 17332 28644
rect 17276 28590 17278 28642
rect 17278 28590 17330 28642
rect 17330 28590 17332 28642
rect 17276 28588 17332 28590
rect 17164 27804 17220 27860
rect 17500 27970 17556 27972
rect 17500 27918 17502 27970
rect 17502 27918 17554 27970
rect 17554 27918 17556 27970
rect 17500 27916 17556 27918
rect 17164 27580 17220 27636
rect 17724 30156 17780 30212
rect 18172 30044 18228 30100
rect 18508 31836 18564 31892
rect 19068 32620 19124 32676
rect 19516 32508 19572 32564
rect 19964 33346 20020 33348
rect 19964 33294 19966 33346
rect 19966 33294 20018 33346
rect 20018 33294 20020 33346
rect 19964 33292 20020 33294
rect 20748 43650 20804 43652
rect 20748 43598 20750 43650
rect 20750 43598 20802 43650
rect 20802 43598 20804 43650
rect 20748 43596 20804 43598
rect 20412 43538 20468 43540
rect 20412 43486 20414 43538
rect 20414 43486 20466 43538
rect 20466 43486 20468 43538
rect 20412 43484 20468 43486
rect 24108 50482 24164 50484
rect 24108 50430 24110 50482
rect 24110 50430 24162 50482
rect 24162 50430 24164 50482
rect 24108 50428 24164 50430
rect 24556 50482 24612 50484
rect 24556 50430 24558 50482
rect 24558 50430 24610 50482
rect 24610 50430 24612 50482
rect 24556 50428 24612 50430
rect 25116 50482 25172 50484
rect 25116 50430 25118 50482
rect 25118 50430 25170 50482
rect 25170 50430 25172 50482
rect 25116 50428 25172 50430
rect 25900 50428 25956 50484
rect 24556 49756 24612 49812
rect 23212 49698 23268 49700
rect 23212 49646 23214 49698
rect 23214 49646 23266 49698
rect 23266 49646 23268 49698
rect 23212 49644 23268 49646
rect 23436 48524 23492 48580
rect 23100 48242 23156 48244
rect 23100 48190 23102 48242
rect 23102 48190 23154 48242
rect 23154 48190 23156 48242
rect 23100 48188 23156 48190
rect 24444 48636 24500 48692
rect 24332 48300 24388 48356
rect 24108 47570 24164 47572
rect 24108 47518 24110 47570
rect 24110 47518 24162 47570
rect 24162 47518 24164 47570
rect 24108 47516 24164 47518
rect 23436 46786 23492 46788
rect 23436 46734 23438 46786
rect 23438 46734 23490 46786
rect 23490 46734 23492 46786
rect 23436 46732 23492 46734
rect 23436 45836 23492 45892
rect 22876 45388 22932 45444
rect 23996 46732 24052 46788
rect 24892 49644 24948 49700
rect 25452 49810 25508 49812
rect 25452 49758 25454 49810
rect 25454 49758 25506 49810
rect 25506 49758 25508 49810
rect 25452 49756 25508 49758
rect 25564 49698 25620 49700
rect 25564 49646 25566 49698
rect 25566 49646 25618 49698
rect 25618 49646 25620 49698
rect 25564 49644 25620 49646
rect 25228 48972 25284 49028
rect 24444 46732 24500 46788
rect 23772 45388 23828 45444
rect 23212 45330 23268 45332
rect 23212 45278 23214 45330
rect 23214 45278 23266 45330
rect 23266 45278 23268 45330
rect 23212 45276 23268 45278
rect 24668 45666 24724 45668
rect 24668 45614 24670 45666
rect 24670 45614 24722 45666
rect 24722 45614 24724 45666
rect 24668 45612 24724 45614
rect 23996 44940 24052 44996
rect 24556 44994 24612 44996
rect 24556 44942 24558 44994
rect 24558 44942 24610 44994
rect 24610 44942 24612 44994
rect 24556 44940 24612 44942
rect 23436 44828 23492 44884
rect 24668 44716 24724 44772
rect 24780 45500 24836 45556
rect 23212 44098 23268 44100
rect 23212 44046 23214 44098
rect 23214 44046 23266 44098
rect 23266 44046 23268 44098
rect 23212 44044 23268 44046
rect 23436 44044 23492 44100
rect 20860 40236 20916 40292
rect 22428 40962 22484 40964
rect 22428 40910 22430 40962
rect 22430 40910 22482 40962
rect 22482 40910 22484 40962
rect 22428 40908 22484 40910
rect 21868 40290 21924 40292
rect 21868 40238 21870 40290
rect 21870 40238 21922 40290
rect 21922 40238 21924 40290
rect 21868 40236 21924 40238
rect 22092 40684 22148 40740
rect 20636 37938 20692 37940
rect 20636 37886 20638 37938
rect 20638 37886 20690 37938
rect 20690 37886 20692 37938
rect 20636 37884 20692 37886
rect 20636 36428 20692 36484
rect 20748 35532 20804 35588
rect 20524 33628 20580 33684
rect 20636 34860 20692 34916
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20300 32956 20356 33012
rect 20412 33516 20468 33572
rect 20044 32900 20100 32902
rect 20748 33964 20804 34020
rect 19852 32562 19908 32564
rect 19852 32510 19854 32562
rect 19854 32510 19906 32562
rect 19906 32510 19908 32562
rect 19852 32508 19908 32510
rect 18508 30940 18564 30996
rect 17836 29260 17892 29316
rect 17836 28642 17892 28644
rect 17836 28590 17838 28642
rect 17838 28590 17890 28642
rect 17890 28590 17892 28642
rect 17836 28588 17892 28590
rect 18396 27916 18452 27972
rect 16940 21644 16996 21700
rect 16492 20076 16548 20132
rect 16716 20636 16772 20692
rect 16156 20018 16212 20020
rect 16156 19966 16158 20018
rect 16158 19966 16210 20018
rect 16210 19966 16212 20018
rect 16156 19964 16212 19966
rect 16604 19740 16660 19796
rect 14700 17500 14756 17556
rect 14812 17724 14868 17780
rect 12460 16044 12516 16100
rect 12684 15874 12740 15876
rect 12684 15822 12686 15874
rect 12686 15822 12738 15874
rect 12738 15822 12740 15874
rect 12684 15820 12740 15822
rect 13132 15426 13188 15428
rect 13132 15374 13134 15426
rect 13134 15374 13186 15426
rect 13186 15374 13188 15426
rect 13132 15372 13188 15374
rect 14364 15372 14420 15428
rect 12012 14530 12068 14532
rect 12012 14478 12014 14530
rect 12014 14478 12066 14530
rect 12066 14478 12068 14530
rect 12012 14476 12068 14478
rect 14028 15148 14084 15204
rect 10220 14306 10276 14308
rect 10220 14254 10222 14306
rect 10222 14254 10274 14306
rect 10274 14254 10276 14306
rect 10220 14252 10276 14254
rect 10668 13468 10724 13524
rect 9548 12236 9604 12292
rect 9212 12124 9268 12180
rect 10108 12178 10164 12180
rect 10108 12126 10110 12178
rect 10110 12126 10162 12178
rect 10162 12126 10164 12178
rect 10108 12124 10164 12126
rect 9324 11282 9380 11284
rect 9324 11230 9326 11282
rect 9326 11230 9378 11282
rect 9378 11230 9380 11282
rect 9324 11228 9380 11230
rect 10332 11954 10388 11956
rect 10332 11902 10334 11954
rect 10334 11902 10386 11954
rect 10386 11902 10388 11954
rect 10332 11900 10388 11902
rect 11676 13692 11732 13748
rect 12124 14252 12180 14308
rect 11564 13468 11620 13524
rect 11004 13020 11060 13076
rect 11900 13074 11956 13076
rect 11900 13022 11902 13074
rect 11902 13022 11954 13074
rect 11954 13022 11956 13074
rect 11900 13020 11956 13022
rect 12124 12908 12180 12964
rect 12348 13746 12404 13748
rect 12348 13694 12350 13746
rect 12350 13694 12402 13746
rect 12402 13694 12404 13746
rect 12348 13692 12404 13694
rect 10668 10668 10724 10724
rect 9884 9212 9940 9268
rect 10892 11228 10948 11284
rect 11676 11228 11732 11284
rect 11004 10892 11060 10948
rect 10892 10834 10948 10836
rect 10892 10782 10894 10834
rect 10894 10782 10946 10834
rect 10946 10782 10948 10834
rect 10892 10780 10948 10782
rect 12124 10892 12180 10948
rect 12012 10834 12068 10836
rect 12012 10782 12014 10834
rect 12014 10782 12066 10834
rect 12066 10782 12068 10834
rect 12012 10780 12068 10782
rect 11452 10444 11508 10500
rect 14364 13692 14420 13748
rect 14588 16882 14644 16884
rect 14588 16830 14590 16882
rect 14590 16830 14642 16882
rect 14642 16830 14644 16882
rect 14588 16828 14644 16830
rect 15708 17778 15764 17780
rect 15708 17726 15710 17778
rect 15710 17726 15762 17778
rect 15762 17726 15764 17778
rect 15708 17724 15764 17726
rect 15148 17554 15204 17556
rect 15148 17502 15150 17554
rect 15150 17502 15202 17554
rect 15202 17502 15204 17554
rect 15148 17500 15204 17502
rect 15036 16268 15092 16324
rect 17724 25564 17780 25620
rect 17612 25394 17668 25396
rect 17612 25342 17614 25394
rect 17614 25342 17666 25394
rect 17666 25342 17668 25394
rect 17612 25340 17668 25342
rect 17500 24946 17556 24948
rect 17500 24894 17502 24946
rect 17502 24894 17554 24946
rect 17554 24894 17556 24946
rect 17500 24892 17556 24894
rect 17724 25228 17780 25284
rect 18396 24332 18452 24388
rect 18060 23884 18116 23940
rect 20300 31554 20356 31556
rect 20300 31502 20302 31554
rect 20302 31502 20354 31554
rect 20354 31502 20356 31554
rect 20300 31500 20356 31502
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 20300 30156 20356 30212
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 18844 29426 18900 29428
rect 18844 29374 18846 29426
rect 18846 29374 18898 29426
rect 18898 29374 18900 29426
rect 18844 29372 18900 29374
rect 19180 28754 19236 28756
rect 19180 28702 19182 28754
rect 19182 28702 19234 28754
rect 19234 28702 19236 28754
rect 19180 28700 19236 28702
rect 19628 28866 19684 28868
rect 19628 28814 19630 28866
rect 19630 28814 19682 28866
rect 19682 28814 19684 28866
rect 19628 28812 19684 28814
rect 19740 28700 19796 28756
rect 18844 28082 18900 28084
rect 18844 28030 18846 28082
rect 18846 28030 18898 28082
rect 18898 28030 18900 28082
rect 18844 28028 18900 28030
rect 19068 27074 19124 27076
rect 19068 27022 19070 27074
rect 19070 27022 19122 27074
rect 19122 27022 19124 27074
rect 19068 27020 19124 27022
rect 19404 27692 19460 27748
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 19964 27970 20020 27972
rect 19964 27918 19966 27970
rect 19966 27918 20018 27970
rect 20018 27918 20020 27970
rect 19964 27916 20020 27918
rect 19628 27692 19684 27748
rect 19516 27468 19572 27524
rect 19292 27356 19348 27412
rect 19964 27074 20020 27076
rect 19964 27022 19966 27074
rect 19966 27022 20018 27074
rect 20018 27022 20020 27074
rect 19964 27020 20020 27022
rect 21644 36482 21700 36484
rect 21644 36430 21646 36482
rect 21646 36430 21698 36482
rect 21698 36430 21700 36482
rect 21644 36428 21700 36430
rect 21868 36316 21924 36372
rect 21532 33292 21588 33348
rect 21644 33234 21700 33236
rect 21644 33182 21646 33234
rect 21646 33182 21698 33234
rect 21698 33182 21700 33234
rect 21644 33180 21700 33182
rect 20860 33068 20916 33124
rect 21644 32284 21700 32340
rect 20412 29932 20468 29988
rect 19404 26962 19460 26964
rect 19404 26910 19406 26962
rect 19406 26910 19458 26962
rect 19458 26910 19460 26962
rect 19404 26908 19460 26910
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19852 25506 19908 25508
rect 19852 25454 19854 25506
rect 19854 25454 19906 25506
rect 19906 25454 19908 25506
rect 19852 25452 19908 25454
rect 19292 24332 19348 24388
rect 18508 20914 18564 20916
rect 18508 20862 18510 20914
rect 18510 20862 18562 20914
rect 18562 20862 18564 20914
rect 18508 20860 18564 20862
rect 18844 20690 18900 20692
rect 18844 20638 18846 20690
rect 18846 20638 18898 20690
rect 18898 20638 18900 20690
rect 18844 20636 18900 20638
rect 19068 20636 19124 20692
rect 17052 19404 17108 19460
rect 16716 16940 16772 16996
rect 15820 16882 15876 16884
rect 15820 16830 15822 16882
rect 15822 16830 15874 16882
rect 15874 16830 15876 16882
rect 15820 16828 15876 16830
rect 17388 16882 17444 16884
rect 17388 16830 17390 16882
rect 17390 16830 17442 16882
rect 17442 16830 17444 16882
rect 17388 16828 17444 16830
rect 18172 17106 18228 17108
rect 18172 17054 18174 17106
rect 18174 17054 18226 17106
rect 18226 17054 18228 17106
rect 18172 17052 18228 17054
rect 16268 16098 16324 16100
rect 16268 16046 16270 16098
rect 16270 16046 16322 16098
rect 16322 16046 16324 16098
rect 16268 16044 16324 16046
rect 15596 15986 15652 15988
rect 15596 15934 15598 15986
rect 15598 15934 15650 15986
rect 15650 15934 15652 15986
rect 15596 15932 15652 15934
rect 15148 15820 15204 15876
rect 16492 16322 16548 16324
rect 16492 16270 16494 16322
rect 16494 16270 16546 16322
rect 16546 16270 16548 16322
rect 16492 16268 16548 16270
rect 16716 16156 16772 16212
rect 17500 16098 17556 16100
rect 17500 16046 17502 16098
rect 17502 16046 17554 16098
rect 17554 16046 17556 16098
rect 17500 16044 17556 16046
rect 18060 16828 18116 16884
rect 17836 16658 17892 16660
rect 17836 16606 17838 16658
rect 17838 16606 17890 16658
rect 17890 16606 17892 16658
rect 17836 16604 17892 16606
rect 16492 15202 16548 15204
rect 16492 15150 16494 15202
rect 16494 15150 16546 15202
rect 16546 15150 16548 15202
rect 16492 15148 16548 15150
rect 14476 13356 14532 13412
rect 14812 13356 14868 13412
rect 13916 12962 13972 12964
rect 13916 12910 13918 12962
rect 13918 12910 13970 12962
rect 13970 12910 13972 12962
rect 13916 12908 13972 12910
rect 14252 12962 14308 12964
rect 14252 12910 14254 12962
rect 14254 12910 14306 12962
rect 14306 12910 14308 12962
rect 14252 12908 14308 12910
rect 12460 12178 12516 12180
rect 12460 12126 12462 12178
rect 12462 12126 12514 12178
rect 12514 12126 12516 12178
rect 12460 12124 12516 12126
rect 13468 12178 13524 12180
rect 13468 12126 13470 12178
rect 13470 12126 13522 12178
rect 13522 12126 13524 12178
rect 13468 12124 13524 12126
rect 12908 12012 12964 12068
rect 12572 11954 12628 11956
rect 12572 11902 12574 11954
rect 12574 11902 12626 11954
rect 12626 11902 12628 11954
rect 12572 11900 12628 11902
rect 13356 11676 13412 11732
rect 12796 11228 12852 11284
rect 13244 10834 13300 10836
rect 13244 10782 13246 10834
rect 13246 10782 13298 10834
rect 13298 10782 13300 10834
rect 13244 10780 13300 10782
rect 12572 10610 12628 10612
rect 12572 10558 12574 10610
rect 12574 10558 12626 10610
rect 12626 10558 12628 10610
rect 12572 10556 12628 10558
rect 13356 10444 13412 10500
rect 11340 9212 11396 9268
rect 14140 12290 14196 12292
rect 14140 12238 14142 12290
rect 14142 12238 14194 12290
rect 14194 12238 14196 12290
rect 14140 12236 14196 12238
rect 14476 12066 14532 12068
rect 14476 12014 14478 12066
rect 14478 12014 14530 12066
rect 14530 12014 14532 12066
rect 14476 12012 14532 12014
rect 14588 11676 14644 11732
rect 14364 11564 14420 11620
rect 14812 12290 14868 12292
rect 14812 12238 14814 12290
rect 14814 12238 14866 12290
rect 14866 12238 14868 12290
rect 14812 12236 14868 12238
rect 15148 12962 15204 12964
rect 15148 12910 15150 12962
rect 15150 12910 15202 12962
rect 15202 12910 15204 12962
rect 15148 12908 15204 12910
rect 15260 11900 15316 11956
rect 15148 11452 15204 11508
rect 14812 11394 14868 11396
rect 14812 11342 14814 11394
rect 14814 11342 14866 11394
rect 14866 11342 14868 11394
rect 14812 11340 14868 11342
rect 16492 15036 16548 15092
rect 16828 15036 16884 15092
rect 16604 14924 16660 14980
rect 16604 14530 16660 14532
rect 16604 14478 16606 14530
rect 16606 14478 16658 14530
rect 16658 14478 16660 14530
rect 16604 14476 16660 14478
rect 15484 13356 15540 13412
rect 16156 13916 16212 13972
rect 17052 15932 17108 15988
rect 17388 15986 17444 15988
rect 17388 15934 17390 15986
rect 17390 15934 17442 15986
rect 17442 15934 17444 15986
rect 17388 15932 17444 15934
rect 16940 14306 16996 14308
rect 16940 14254 16942 14306
rect 16942 14254 16994 14306
rect 16994 14254 16996 14306
rect 16940 14252 16996 14254
rect 16380 13858 16436 13860
rect 16380 13806 16382 13858
rect 16382 13806 16434 13858
rect 16434 13806 16436 13858
rect 16380 13804 16436 13806
rect 17276 14530 17332 14532
rect 17276 14478 17278 14530
rect 17278 14478 17330 14530
rect 17330 14478 17332 14530
rect 17276 14476 17332 14478
rect 17164 14252 17220 14308
rect 17052 13804 17108 13860
rect 17612 13804 17668 13860
rect 17724 13916 17780 13972
rect 15932 13746 15988 13748
rect 15932 13694 15934 13746
rect 15934 13694 15986 13746
rect 15986 13694 15988 13746
rect 15932 13692 15988 13694
rect 18620 16716 18676 16772
rect 18508 16604 18564 16660
rect 18172 16210 18228 16212
rect 18172 16158 18174 16210
rect 18174 16158 18226 16210
rect 18226 16158 18228 16210
rect 18172 16156 18228 16158
rect 18620 15426 18676 15428
rect 18620 15374 18622 15426
rect 18622 15374 18674 15426
rect 18674 15374 18676 15426
rect 18620 15372 18676 15374
rect 18844 15202 18900 15204
rect 18844 15150 18846 15202
rect 18846 15150 18898 15202
rect 18898 15150 18900 15202
rect 18844 15148 18900 15150
rect 18284 13858 18340 13860
rect 18284 13806 18286 13858
rect 18286 13806 18338 13858
rect 18338 13806 18340 13858
rect 18284 13804 18340 13806
rect 18396 14476 18452 14532
rect 18844 14252 18900 14308
rect 18508 13746 18564 13748
rect 18508 13694 18510 13746
rect 18510 13694 18562 13746
rect 18562 13694 18564 13746
rect 18508 13692 18564 13694
rect 18732 13634 18788 13636
rect 18732 13582 18734 13634
rect 18734 13582 18786 13634
rect 18786 13582 18788 13634
rect 18732 13580 18788 13582
rect 18844 13468 18900 13524
rect 19068 14530 19124 14532
rect 19068 14478 19070 14530
rect 19070 14478 19122 14530
rect 19122 14478 19124 14530
rect 19068 14476 19124 14478
rect 19068 13580 19124 13636
rect 15932 11564 15988 11620
rect 14028 11282 14084 11284
rect 14028 11230 14030 11282
rect 14030 11230 14082 11282
rect 14082 11230 14084 11282
rect 14028 11228 14084 11230
rect 15148 11282 15204 11284
rect 15148 11230 15150 11282
rect 15150 11230 15202 11282
rect 15202 11230 15204 11282
rect 15148 11228 15204 11230
rect 13916 10556 13972 10612
rect 13692 9548 13748 9604
rect 11340 8428 11396 8484
rect 9548 8034 9604 8036
rect 9548 7982 9550 8034
rect 9550 7982 9602 8034
rect 9602 7982 9604 8034
rect 9548 7980 9604 7982
rect 10780 7980 10836 8036
rect 8988 7698 9044 7700
rect 8988 7646 8990 7698
rect 8990 7646 9042 7698
rect 9042 7646 9044 7698
rect 8988 7644 9044 7646
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 3724 4226 3780 4228
rect 3724 4174 3726 4226
rect 3726 4174 3778 4226
rect 3778 4174 3780 4226
rect 3724 4172 3780 4174
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 13356 8428 13412 8484
rect 12124 7532 12180 7588
rect 14364 11116 14420 11172
rect 15260 11170 15316 11172
rect 15260 11118 15262 11170
rect 15262 11118 15314 11170
rect 15314 11118 15316 11170
rect 15260 11116 15316 11118
rect 15820 11394 15876 11396
rect 15820 11342 15822 11394
rect 15822 11342 15874 11394
rect 15874 11342 15876 11394
rect 15820 11340 15876 11342
rect 16604 11452 16660 11508
rect 19292 17052 19348 17108
rect 19740 25282 19796 25284
rect 19740 25230 19742 25282
rect 19742 25230 19794 25282
rect 19794 25230 19796 25282
rect 19740 25228 19796 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19852 24722 19908 24724
rect 19852 24670 19854 24722
rect 19854 24670 19906 24722
rect 19906 24670 19908 24722
rect 19852 24668 19908 24670
rect 20300 29484 20356 29540
rect 20412 29036 20468 29092
rect 20636 30098 20692 30100
rect 20636 30046 20638 30098
rect 20638 30046 20690 30098
rect 20690 30046 20692 30098
rect 20636 30044 20692 30046
rect 21420 29986 21476 29988
rect 21420 29934 21422 29986
rect 21422 29934 21474 29986
rect 21474 29934 21476 29986
rect 21420 29932 21476 29934
rect 21420 29036 21476 29092
rect 20524 28028 20580 28084
rect 20300 26908 20356 26964
rect 20300 25282 20356 25284
rect 20300 25230 20302 25282
rect 20302 25230 20354 25282
rect 20354 25230 20356 25282
rect 20300 25228 20356 25230
rect 20524 25116 20580 25172
rect 20300 24722 20356 24724
rect 20300 24670 20302 24722
rect 20302 24670 20354 24722
rect 20354 24670 20356 24722
rect 20300 24668 20356 24670
rect 20076 23660 20132 23716
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20412 22092 20468 22148
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 19628 20690 19684 20692
rect 19628 20638 19630 20690
rect 19630 20638 19682 20690
rect 19682 20638 19684 20690
rect 19628 20636 19684 20638
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19628 16716 19684 16772
rect 21868 30210 21924 30212
rect 21868 30158 21870 30210
rect 21870 30158 21922 30210
rect 21922 30158 21924 30210
rect 21868 30156 21924 30158
rect 21980 30828 22036 30884
rect 21756 28700 21812 28756
rect 21980 28364 22036 28420
rect 21980 27916 22036 27972
rect 21084 25116 21140 25172
rect 20636 24834 20692 24836
rect 20636 24782 20638 24834
rect 20638 24782 20690 24834
rect 20690 24782 20692 24834
rect 20636 24780 20692 24782
rect 20636 23436 20692 23492
rect 21420 23660 21476 23716
rect 20636 22876 20692 22932
rect 21868 24946 21924 24948
rect 21868 24894 21870 24946
rect 21870 24894 21922 24946
rect 21922 24894 21924 24946
rect 21868 24892 21924 24894
rect 22652 40684 22708 40740
rect 22316 40572 22372 40628
rect 22988 41970 23044 41972
rect 22988 41918 22990 41970
rect 22990 41918 23042 41970
rect 23042 41918 23044 41970
rect 22988 41916 23044 41918
rect 23436 41916 23492 41972
rect 22988 41244 23044 41300
rect 23436 41692 23492 41748
rect 23436 40684 23492 40740
rect 23324 40626 23380 40628
rect 23324 40574 23326 40626
rect 23326 40574 23378 40626
rect 23378 40574 23380 40626
rect 23324 40572 23380 40574
rect 23324 40402 23380 40404
rect 23324 40350 23326 40402
rect 23326 40350 23378 40402
rect 23378 40350 23380 40402
rect 23324 40348 23380 40350
rect 23884 42028 23940 42084
rect 23772 41970 23828 41972
rect 23772 41918 23774 41970
rect 23774 41918 23826 41970
rect 23826 41918 23828 41970
rect 23772 41916 23828 41918
rect 23660 41132 23716 41188
rect 23996 41468 24052 41524
rect 23996 40908 24052 40964
rect 24220 41244 24276 41300
rect 24668 41804 24724 41860
rect 24556 40402 24612 40404
rect 24556 40350 24558 40402
rect 24558 40350 24610 40402
rect 24610 40350 24612 40402
rect 24556 40348 24612 40350
rect 25004 48524 25060 48580
rect 25228 48242 25284 48244
rect 25228 48190 25230 48242
rect 25230 48190 25282 48242
rect 25282 48190 25284 48242
rect 25228 48188 25284 48190
rect 25676 48636 25732 48692
rect 27692 50594 27748 50596
rect 27692 50542 27694 50594
rect 27694 50542 27746 50594
rect 27746 50542 27748 50594
rect 27692 50540 27748 50542
rect 27356 50482 27412 50484
rect 27356 50430 27358 50482
rect 27358 50430 27410 50482
rect 27410 50430 27412 50482
rect 27356 50428 27412 50430
rect 27244 49308 27300 49364
rect 27356 49420 27412 49476
rect 26684 48972 26740 49028
rect 27020 48972 27076 49028
rect 26572 48412 26628 48468
rect 25564 48354 25620 48356
rect 25564 48302 25566 48354
rect 25566 48302 25618 48354
rect 25618 48302 25620 48354
rect 25564 48300 25620 48302
rect 26236 48242 26292 48244
rect 26236 48190 26238 48242
rect 26238 48190 26290 48242
rect 26290 48190 26292 48242
rect 26236 48188 26292 48190
rect 27132 48636 27188 48692
rect 27132 48466 27188 48468
rect 27132 48414 27134 48466
rect 27134 48414 27186 48466
rect 27186 48414 27188 48466
rect 27132 48412 27188 48414
rect 26012 47516 26068 47572
rect 26348 47458 26404 47460
rect 26348 47406 26350 47458
rect 26350 47406 26402 47458
rect 26402 47406 26404 47458
rect 26348 47404 26404 47406
rect 25452 47346 25508 47348
rect 25452 47294 25454 47346
rect 25454 47294 25506 47346
rect 25506 47294 25508 47346
rect 25452 47292 25508 47294
rect 26572 47292 26628 47348
rect 26908 48300 26964 48356
rect 26236 47234 26292 47236
rect 26236 47182 26238 47234
rect 26238 47182 26290 47234
rect 26290 47182 26292 47234
rect 26236 47180 26292 47182
rect 25452 45666 25508 45668
rect 25452 45614 25454 45666
rect 25454 45614 25506 45666
rect 25506 45614 25508 45666
rect 25452 45612 25508 45614
rect 25228 45276 25284 45332
rect 25228 44268 25284 44324
rect 25564 44268 25620 44324
rect 25116 43708 25172 43764
rect 25900 43538 25956 43540
rect 25900 43486 25902 43538
rect 25902 43486 25954 43538
rect 25954 43486 25956 43538
rect 25900 43484 25956 43486
rect 26236 44098 26292 44100
rect 26236 44046 26238 44098
rect 26238 44046 26290 44098
rect 26290 44046 26292 44098
rect 26236 44044 26292 44046
rect 27020 47516 27076 47572
rect 27132 47180 27188 47236
rect 27244 46844 27300 46900
rect 27580 48242 27636 48244
rect 27580 48190 27582 48242
rect 27582 48190 27634 48242
rect 27634 48190 27636 48242
rect 27580 48188 27636 48190
rect 28588 50428 28644 50484
rect 27916 48748 27972 48804
rect 28476 49420 28532 49476
rect 28252 47458 28308 47460
rect 28252 47406 28254 47458
rect 28254 47406 28306 47458
rect 28306 47406 28308 47458
rect 28252 47404 28308 47406
rect 27468 46898 27524 46900
rect 27468 46846 27470 46898
rect 27470 46846 27522 46898
rect 27522 46846 27524 46898
rect 27468 46844 27524 46846
rect 26012 43260 26068 43316
rect 26124 41970 26180 41972
rect 26124 41918 26126 41970
rect 26126 41918 26178 41970
rect 26178 41918 26180 41970
rect 26124 41916 26180 41918
rect 27020 44098 27076 44100
rect 27020 44046 27022 44098
rect 27022 44046 27074 44098
rect 27074 44046 27076 44098
rect 27020 44044 27076 44046
rect 28140 47346 28196 47348
rect 28140 47294 28142 47346
rect 28142 47294 28194 47346
rect 28194 47294 28196 47346
rect 28140 47292 28196 47294
rect 30716 49420 30772 49476
rect 28476 46620 28532 46676
rect 27468 43708 27524 43764
rect 28364 44940 28420 44996
rect 28364 44604 28420 44660
rect 27132 43538 27188 43540
rect 27132 43486 27134 43538
rect 27134 43486 27186 43538
rect 27186 43486 27188 43538
rect 27132 43484 27188 43486
rect 27244 43426 27300 43428
rect 27244 43374 27246 43426
rect 27246 43374 27298 43426
rect 27298 43374 27300 43426
rect 27244 43372 27300 43374
rect 29148 48748 29204 48804
rect 30940 48802 30996 48804
rect 30940 48750 30942 48802
rect 30942 48750 30994 48802
rect 30994 48750 30996 48802
rect 30940 48748 30996 48750
rect 31052 48636 31108 48692
rect 29932 47346 29988 47348
rect 29932 47294 29934 47346
rect 29934 47294 29986 47346
rect 29986 47294 29988 47346
rect 29932 47292 29988 47294
rect 31724 49698 31780 49700
rect 31724 49646 31726 49698
rect 31726 49646 31778 49698
rect 31778 49646 31780 49698
rect 31724 49644 31780 49646
rect 32060 49084 32116 49140
rect 35196 49418 35252 49420
rect 35196 49366 35198 49418
rect 35198 49366 35250 49418
rect 35250 49366 35252 49418
rect 35196 49364 35252 49366
rect 35300 49418 35356 49420
rect 35300 49366 35302 49418
rect 35302 49366 35354 49418
rect 35354 49366 35356 49418
rect 35300 49364 35356 49366
rect 35404 49418 35460 49420
rect 35404 49366 35406 49418
rect 35406 49366 35458 49418
rect 35458 49366 35460 49418
rect 35404 49364 35460 49366
rect 35644 49420 35700 49476
rect 35196 49084 35252 49140
rect 36764 48860 36820 48916
rect 33964 48748 34020 48804
rect 35532 48748 35588 48804
rect 32284 48636 32340 48692
rect 31612 48130 31668 48132
rect 31612 48078 31614 48130
rect 31614 48078 31666 48130
rect 31666 48078 31668 48130
rect 31612 48076 31668 48078
rect 31948 48018 32004 48020
rect 31948 47966 31950 48018
rect 31950 47966 32002 48018
rect 32002 47966 32004 48018
rect 31948 47964 32004 47966
rect 29932 46562 29988 46564
rect 29932 46510 29934 46562
rect 29934 46510 29986 46562
rect 29986 46510 29988 46562
rect 29932 46508 29988 46510
rect 30268 46620 30324 46676
rect 30940 46844 30996 46900
rect 32060 46844 32116 46900
rect 33180 47964 33236 48020
rect 35196 47850 35252 47852
rect 35196 47798 35198 47850
rect 35198 47798 35250 47850
rect 35250 47798 35252 47850
rect 35196 47796 35252 47798
rect 35300 47850 35356 47852
rect 35300 47798 35302 47850
rect 35302 47798 35354 47850
rect 35354 47798 35356 47850
rect 35300 47796 35356 47798
rect 35404 47850 35460 47852
rect 35404 47798 35406 47850
rect 35406 47798 35458 47850
rect 35458 47798 35460 47850
rect 35404 47796 35460 47798
rect 33740 47516 33796 47572
rect 27356 43260 27412 43316
rect 28588 43484 28644 43540
rect 28588 43260 28644 43316
rect 26348 41468 26404 41524
rect 27356 41804 27412 41860
rect 26796 41410 26852 41412
rect 26796 41358 26798 41410
rect 26798 41358 26850 41410
rect 26850 41358 26852 41410
rect 26796 41356 26852 41358
rect 26012 41244 26068 41300
rect 26572 41186 26628 41188
rect 26572 41134 26574 41186
rect 26574 41134 26626 41186
rect 26626 41134 26628 41186
rect 26572 41132 26628 41134
rect 25452 40460 25508 40516
rect 27916 41244 27972 41300
rect 25900 40402 25956 40404
rect 25900 40350 25902 40402
rect 25902 40350 25954 40402
rect 25954 40350 25956 40402
rect 25900 40348 25956 40350
rect 24444 37996 24500 38052
rect 25340 37324 25396 37380
rect 25788 38050 25844 38052
rect 25788 37998 25790 38050
rect 25790 37998 25842 38050
rect 25842 37998 25844 38050
rect 25788 37996 25844 37998
rect 26348 38050 26404 38052
rect 26348 37998 26350 38050
rect 26350 37998 26402 38050
rect 26402 37998 26404 38050
rect 26348 37996 26404 37998
rect 26908 37996 26964 38052
rect 26460 37548 26516 37604
rect 26796 37378 26852 37380
rect 26796 37326 26798 37378
rect 26798 37326 26850 37378
rect 26850 37326 26852 37378
rect 26796 37324 26852 37326
rect 26236 37266 26292 37268
rect 26236 37214 26238 37266
rect 26238 37214 26290 37266
rect 26290 37214 26292 37266
rect 26236 37212 26292 37214
rect 22876 36876 22932 36932
rect 22316 36316 22372 36372
rect 24668 36316 24724 36372
rect 22204 34860 22260 34916
rect 24556 34914 24612 34916
rect 24556 34862 24558 34914
rect 24558 34862 24610 34914
rect 24610 34862 24612 34914
rect 24556 34860 24612 34862
rect 24220 34690 24276 34692
rect 24220 34638 24222 34690
rect 24222 34638 24274 34690
rect 24274 34638 24276 34690
rect 24220 34636 24276 34638
rect 24892 34690 24948 34692
rect 24892 34638 24894 34690
rect 24894 34638 24946 34690
rect 24946 34638 24948 34690
rect 24892 34636 24948 34638
rect 24668 34524 24724 34580
rect 23772 34076 23828 34132
rect 23324 34018 23380 34020
rect 23324 33966 23326 34018
rect 23326 33966 23378 34018
rect 23378 33966 23380 34018
rect 23324 33964 23380 33966
rect 23996 33964 24052 34020
rect 22764 33180 22820 33236
rect 23436 33122 23492 33124
rect 23436 33070 23438 33122
rect 23438 33070 23490 33122
rect 23490 33070 23492 33122
rect 23436 33068 23492 33070
rect 22988 32508 23044 32564
rect 23548 32562 23604 32564
rect 23548 32510 23550 32562
rect 23550 32510 23602 32562
rect 23602 32510 23604 32562
rect 23548 32508 23604 32510
rect 23436 31836 23492 31892
rect 22540 30044 22596 30100
rect 22428 29820 22484 29876
rect 22204 28082 22260 28084
rect 22204 28030 22206 28082
rect 22206 28030 22258 28082
rect 22258 28030 22260 28082
rect 22204 28028 22260 28030
rect 24780 33964 24836 34020
rect 24108 33122 24164 33124
rect 24108 33070 24110 33122
rect 24110 33070 24162 33122
rect 24162 33070 24164 33122
rect 24108 33068 24164 33070
rect 24108 32620 24164 32676
rect 23660 31666 23716 31668
rect 23660 31614 23662 31666
rect 23662 31614 23714 31666
rect 23714 31614 23716 31666
rect 23660 31612 23716 31614
rect 23884 30380 23940 30436
rect 24332 31388 24388 31444
rect 24220 31052 24276 31108
rect 24444 31276 24500 31332
rect 23324 30098 23380 30100
rect 23324 30046 23326 30098
rect 23326 30046 23378 30098
rect 23378 30046 23380 30098
rect 23324 30044 23380 30046
rect 23212 29650 23268 29652
rect 23212 29598 23214 29650
rect 23214 29598 23266 29650
rect 23266 29598 23268 29650
rect 23212 29596 23268 29598
rect 22876 29538 22932 29540
rect 22876 29486 22878 29538
rect 22878 29486 22930 29538
rect 22930 29486 22932 29538
rect 22876 29484 22932 29486
rect 23436 28476 23492 28532
rect 22428 27580 22484 27636
rect 22204 27468 22260 27524
rect 22540 27468 22596 27524
rect 22204 27020 22260 27076
rect 22316 24946 22372 24948
rect 22316 24894 22318 24946
rect 22318 24894 22370 24946
rect 22370 24894 22372 24946
rect 22316 24892 22372 24894
rect 22092 23436 22148 23492
rect 21756 22316 21812 22372
rect 21868 21810 21924 21812
rect 21868 21758 21870 21810
rect 21870 21758 21922 21810
rect 21922 21758 21924 21810
rect 21868 21756 21924 21758
rect 22204 21756 22260 21812
rect 21532 21308 21588 21364
rect 22652 21810 22708 21812
rect 22652 21758 22654 21810
rect 22654 21758 22706 21810
rect 22706 21758 22708 21810
rect 22652 21756 22708 21758
rect 22316 21308 22372 21364
rect 20972 20188 21028 20244
rect 21532 18956 21588 19012
rect 22204 20188 22260 20244
rect 22092 19628 22148 19684
rect 22092 17724 22148 17780
rect 23436 27858 23492 27860
rect 23436 27806 23438 27858
rect 23438 27806 23490 27858
rect 23490 27806 23492 27858
rect 23436 27804 23492 27806
rect 23772 29986 23828 29988
rect 23772 29934 23774 29986
rect 23774 29934 23826 29986
rect 23826 29934 23828 29986
rect 23772 29932 23828 29934
rect 23996 28476 24052 28532
rect 23996 28082 24052 28084
rect 23996 28030 23998 28082
rect 23998 28030 24050 28082
rect 24050 28030 24052 28082
rect 23996 28028 24052 28030
rect 23772 27916 23828 27972
rect 23548 26796 23604 26852
rect 22988 25228 23044 25284
rect 22988 24834 23044 24836
rect 22988 24782 22990 24834
rect 22990 24782 23042 24834
rect 23042 24782 23044 24834
rect 22988 24780 23044 24782
rect 22988 21644 23044 21700
rect 23212 21586 23268 21588
rect 23212 21534 23214 21586
rect 23214 21534 23266 21586
rect 23266 21534 23268 21586
rect 23212 21532 23268 21534
rect 23660 22316 23716 22372
rect 23548 21756 23604 21812
rect 23436 19628 23492 19684
rect 21868 17666 21924 17668
rect 21868 17614 21870 17666
rect 21870 17614 21922 17666
rect 21922 17614 21924 17666
rect 21868 17612 21924 17614
rect 20524 16156 20580 16212
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19292 15372 19348 15428
rect 19740 15426 19796 15428
rect 19740 15374 19742 15426
rect 19742 15374 19794 15426
rect 19794 15374 19796 15426
rect 19740 15372 19796 15374
rect 21532 16716 21588 16772
rect 20636 14476 20692 14532
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 19516 13634 19572 13636
rect 19516 13582 19518 13634
rect 19518 13582 19570 13634
rect 19570 13582 19572 13634
rect 19516 13580 19572 13582
rect 19404 13522 19460 13524
rect 19404 13470 19406 13522
rect 19406 13470 19458 13522
rect 19458 13470 19460 13522
rect 19404 13468 19460 13470
rect 18844 11340 18900 11396
rect 15484 9548 15540 9604
rect 16716 9602 16772 9604
rect 16716 9550 16718 9602
rect 16718 9550 16770 9602
rect 16770 9550 16772 9602
rect 16716 9548 16772 9550
rect 20300 13746 20356 13748
rect 20300 13694 20302 13746
rect 20302 13694 20354 13746
rect 20354 13694 20356 13746
rect 20300 13692 20356 13694
rect 21644 16604 21700 16660
rect 22540 19010 22596 19012
rect 22540 18958 22542 19010
rect 22542 18958 22594 19010
rect 22594 18958 22596 19010
rect 22540 18956 22596 18958
rect 22876 18508 22932 18564
rect 22876 17612 22932 17668
rect 22316 16770 22372 16772
rect 22316 16718 22318 16770
rect 22318 16718 22370 16770
rect 22370 16718 22372 16770
rect 22316 16716 22372 16718
rect 22204 16604 22260 16660
rect 22652 16604 22708 16660
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 20748 12124 20804 12180
rect 19180 11954 19236 11956
rect 19180 11902 19182 11954
rect 19182 11902 19234 11954
rect 19234 11902 19236 11954
rect 19180 11900 19236 11902
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19068 10780 19124 10836
rect 21420 11676 21476 11732
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 16828 8428 16884 8484
rect 20300 8930 20356 8932
rect 20300 8878 20302 8930
rect 20302 8878 20354 8930
rect 20354 8878 20356 8930
rect 20300 8876 20356 8878
rect 18172 8316 18228 8372
rect 19404 8370 19460 8372
rect 19404 8318 19406 8370
rect 19406 8318 19458 8370
rect 19458 8318 19460 8370
rect 19404 8316 19460 8318
rect 19628 8204 19684 8260
rect 19516 7644 19572 7700
rect 14140 7532 14196 7588
rect 18284 7532 18340 7588
rect 13580 6636 13636 6692
rect 16156 6748 16212 6804
rect 14700 6636 14756 6692
rect 15036 6690 15092 6692
rect 15036 6638 15038 6690
rect 15038 6638 15090 6690
rect 15090 6638 15092 6690
rect 15036 6636 15092 6638
rect 15372 6690 15428 6692
rect 15372 6638 15374 6690
rect 15374 6638 15426 6690
rect 15426 6638 15428 6690
rect 15372 6636 15428 6638
rect 20188 8428 20244 8484
rect 19740 8146 19796 8148
rect 19740 8094 19742 8146
rect 19742 8094 19794 8146
rect 19794 8094 19796 8146
rect 19740 8092 19796 8094
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 23212 16604 23268 16660
rect 23660 18508 23716 18564
rect 23660 17554 23716 17556
rect 23660 17502 23662 17554
rect 23662 17502 23714 17554
rect 23714 17502 23716 17554
rect 23660 17500 23716 17502
rect 23548 16716 23604 16772
rect 21868 13468 21924 13524
rect 22876 13468 22932 13524
rect 22428 12796 22484 12852
rect 21868 12178 21924 12180
rect 21868 12126 21870 12178
rect 21870 12126 21922 12178
rect 21922 12126 21924 12178
rect 21868 12124 21924 12126
rect 21532 11116 21588 11172
rect 22316 12178 22372 12180
rect 22316 12126 22318 12178
rect 22318 12126 22370 12178
rect 22370 12126 22372 12178
rect 22316 12124 22372 12126
rect 22204 11676 22260 11732
rect 21308 9884 21364 9940
rect 22092 9884 22148 9940
rect 22764 9884 22820 9940
rect 24108 26796 24164 26852
rect 23884 25506 23940 25508
rect 23884 25454 23886 25506
rect 23886 25454 23938 25506
rect 23938 25454 23940 25506
rect 23884 25452 23940 25454
rect 24220 27692 24276 27748
rect 24108 25340 24164 25396
rect 24332 22316 24388 22372
rect 23996 22146 24052 22148
rect 23996 22094 23998 22146
rect 23998 22094 24050 22146
rect 24050 22094 24052 22146
rect 23996 22092 24052 22094
rect 23884 21698 23940 21700
rect 23884 21646 23886 21698
rect 23886 21646 23938 21698
rect 23938 21646 23940 21698
rect 23884 21644 23940 21646
rect 23996 19852 24052 19908
rect 24556 31052 24612 31108
rect 24668 30994 24724 30996
rect 24668 30942 24670 30994
rect 24670 30942 24722 30994
rect 24722 30942 24724 30994
rect 24668 30940 24724 30942
rect 24556 29986 24612 29988
rect 24556 29934 24558 29986
rect 24558 29934 24610 29986
rect 24610 29934 24612 29986
rect 24556 29932 24612 29934
rect 24668 27244 24724 27300
rect 24556 25506 24612 25508
rect 24556 25454 24558 25506
rect 24558 25454 24610 25506
rect 24610 25454 24612 25506
rect 24556 25452 24612 25454
rect 24668 24946 24724 24948
rect 24668 24894 24670 24946
rect 24670 24894 24722 24946
rect 24722 24894 24724 24946
rect 24668 24892 24724 24894
rect 24668 21868 24724 21924
rect 26908 36876 26964 36932
rect 25452 34636 25508 34692
rect 26012 33964 26068 34020
rect 25452 32732 25508 32788
rect 25340 32060 25396 32116
rect 25452 31948 25508 32004
rect 25004 31276 25060 31332
rect 25116 31052 25172 31108
rect 25228 30994 25284 30996
rect 25228 30942 25230 30994
rect 25230 30942 25282 30994
rect 25282 30942 25284 30994
rect 25228 30940 25284 30942
rect 25340 29820 25396 29876
rect 25452 31500 25508 31556
rect 25228 29596 25284 29652
rect 25116 28924 25172 28980
rect 24892 28642 24948 28644
rect 24892 28590 24894 28642
rect 24894 28590 24946 28642
rect 24946 28590 24948 28642
rect 24892 28588 24948 28590
rect 25004 27074 25060 27076
rect 25004 27022 25006 27074
rect 25006 27022 25058 27074
rect 25058 27022 25060 27074
rect 25004 27020 25060 27022
rect 25340 28588 25396 28644
rect 25228 26962 25284 26964
rect 25228 26910 25230 26962
rect 25230 26910 25282 26962
rect 25282 26910 25284 26962
rect 25228 26908 25284 26910
rect 25340 26796 25396 26852
rect 26236 32786 26292 32788
rect 26236 32734 26238 32786
rect 26238 32734 26290 32786
rect 26290 32734 26292 32786
rect 26236 32732 26292 32734
rect 26236 31948 26292 32004
rect 25788 31612 25844 31668
rect 25788 30828 25844 30884
rect 25564 30210 25620 30212
rect 25564 30158 25566 30210
rect 25566 30158 25618 30210
rect 25618 30158 25620 30210
rect 25564 30156 25620 30158
rect 26236 30210 26292 30212
rect 26236 30158 26238 30210
rect 26238 30158 26290 30210
rect 26290 30158 26292 30210
rect 26236 30156 26292 30158
rect 26124 29314 26180 29316
rect 26124 29262 26126 29314
rect 26126 29262 26178 29314
rect 26178 29262 26180 29314
rect 26124 29260 26180 29262
rect 25788 28754 25844 28756
rect 25788 28702 25790 28754
rect 25790 28702 25842 28754
rect 25842 28702 25844 28754
rect 25788 28700 25844 28702
rect 26236 28700 26292 28756
rect 25564 28588 25620 28644
rect 25452 27916 25508 27972
rect 25228 25394 25284 25396
rect 25228 25342 25230 25394
rect 25230 25342 25282 25394
rect 25282 25342 25284 25394
rect 25228 25340 25284 25342
rect 25228 23714 25284 23716
rect 25228 23662 25230 23714
rect 25230 23662 25282 23714
rect 25282 23662 25284 23714
rect 25228 23660 25284 23662
rect 24780 21532 24836 21588
rect 24780 20130 24836 20132
rect 24780 20078 24782 20130
rect 24782 20078 24834 20130
rect 24834 20078 24836 20130
rect 24780 20076 24836 20078
rect 25340 19906 25396 19908
rect 25340 19854 25342 19906
rect 25342 19854 25394 19906
rect 25394 19854 25396 19906
rect 25340 19852 25396 19854
rect 25676 28364 25732 28420
rect 25676 27020 25732 27076
rect 25788 26796 25844 26852
rect 26236 26460 26292 26516
rect 26460 30882 26516 30884
rect 26460 30830 26462 30882
rect 26462 30830 26514 30882
rect 26514 30830 26516 30882
rect 26460 30828 26516 30830
rect 26460 29260 26516 29316
rect 26460 28924 26516 28980
rect 26460 28588 26516 28644
rect 26460 26908 26516 26964
rect 25564 24892 25620 24948
rect 25788 25452 25844 25508
rect 25788 24946 25844 24948
rect 25788 24894 25790 24946
rect 25790 24894 25842 24946
rect 25842 24894 25844 24946
rect 25788 24892 25844 24894
rect 25676 23436 25732 23492
rect 25900 22146 25956 22148
rect 25900 22094 25902 22146
rect 25902 22094 25954 22146
rect 25954 22094 25956 22146
rect 25900 22092 25956 22094
rect 25564 21868 25620 21924
rect 25788 20130 25844 20132
rect 25788 20078 25790 20130
rect 25790 20078 25842 20130
rect 25842 20078 25844 20130
rect 25788 20076 25844 20078
rect 25564 20018 25620 20020
rect 25564 19966 25566 20018
rect 25566 19966 25618 20018
rect 25618 19966 25620 20018
rect 25564 19964 25620 19966
rect 26348 25618 26404 25620
rect 26348 25566 26350 25618
rect 26350 25566 26402 25618
rect 26402 25566 26404 25618
rect 26348 25564 26404 25566
rect 26236 24668 26292 24724
rect 26124 24050 26180 24052
rect 26124 23998 26126 24050
rect 26126 23998 26178 24050
rect 26178 23998 26180 24050
rect 26124 23996 26180 23998
rect 26124 23660 26180 23716
rect 25340 18562 25396 18564
rect 25340 18510 25342 18562
rect 25342 18510 25394 18562
rect 25394 18510 25396 18562
rect 25340 18508 25396 18510
rect 26012 18508 26068 18564
rect 26908 28754 26964 28756
rect 26908 28702 26910 28754
rect 26910 28702 26962 28754
rect 26962 28702 26964 28754
rect 26908 28700 26964 28702
rect 27132 34188 27188 34244
rect 27356 29820 27412 29876
rect 27356 28754 27412 28756
rect 27356 28702 27358 28754
rect 27358 28702 27410 28754
rect 27410 28702 27412 28754
rect 27356 28700 27412 28702
rect 28588 40684 28644 40740
rect 30156 45388 30212 45444
rect 29260 43538 29316 43540
rect 29260 43486 29262 43538
rect 29262 43486 29314 43538
rect 29314 43486 29316 43538
rect 29260 43484 29316 43486
rect 29708 43372 29764 43428
rect 29372 43314 29428 43316
rect 29372 43262 29374 43314
rect 29374 43262 29426 43314
rect 29426 43262 29428 43314
rect 29372 43260 29428 43262
rect 30044 42364 30100 42420
rect 29148 41244 29204 41300
rect 29148 40402 29204 40404
rect 29148 40350 29150 40402
rect 29150 40350 29202 40402
rect 29202 40350 29204 40402
rect 29148 40348 29204 40350
rect 30940 45388 30996 45444
rect 32284 45276 32340 45332
rect 31500 44994 31556 44996
rect 31500 44942 31502 44994
rect 31502 44942 31554 44994
rect 31554 44942 31556 44994
rect 31500 44940 31556 44942
rect 32060 44434 32116 44436
rect 32060 44382 32062 44434
rect 32062 44382 32114 44434
rect 32114 44382 32116 44434
rect 32060 44380 32116 44382
rect 33516 46786 33572 46788
rect 33516 46734 33518 46786
rect 33518 46734 33570 46786
rect 33570 46734 33572 46786
rect 33516 46732 33572 46734
rect 35308 47570 35364 47572
rect 35308 47518 35310 47570
rect 35310 47518 35362 47570
rect 35362 47518 35364 47570
rect 35308 47516 35364 47518
rect 37436 49810 37492 49812
rect 37436 49758 37438 49810
rect 37438 49758 37490 49810
rect 37490 49758 37492 49810
rect 37436 49756 37492 49758
rect 36876 48748 36932 48804
rect 37100 47516 37156 47572
rect 37212 48860 37268 48916
rect 36204 46562 36260 46564
rect 36204 46510 36206 46562
rect 36206 46510 36258 46562
rect 36258 46510 36260 46562
rect 36204 46508 36260 46510
rect 37100 46508 37156 46564
rect 35196 46282 35252 46284
rect 35196 46230 35198 46282
rect 35198 46230 35250 46282
rect 35250 46230 35252 46282
rect 35196 46228 35252 46230
rect 35300 46282 35356 46284
rect 35300 46230 35302 46282
rect 35302 46230 35354 46282
rect 35354 46230 35356 46282
rect 35300 46228 35356 46230
rect 35404 46282 35460 46284
rect 35404 46230 35406 46282
rect 35406 46230 35458 46282
rect 35458 46230 35460 46282
rect 35404 46228 35460 46230
rect 32844 44940 32900 44996
rect 33292 44882 33348 44884
rect 33292 44830 33294 44882
rect 33294 44830 33346 44882
rect 33346 44830 33348 44882
rect 33292 44828 33348 44830
rect 32844 44434 32900 44436
rect 32844 44382 32846 44434
rect 32846 44382 32898 44434
rect 32898 44382 32900 44434
rect 32844 44380 32900 44382
rect 33404 44380 33460 44436
rect 30492 42364 30548 42420
rect 32732 42530 32788 42532
rect 32732 42478 32734 42530
rect 32734 42478 32786 42530
rect 32786 42478 32788 42530
rect 32732 42476 32788 42478
rect 31948 41858 32004 41860
rect 31948 41806 31950 41858
rect 31950 41806 32002 41858
rect 32002 41806 32004 41858
rect 31948 41804 32004 41806
rect 33292 42476 33348 42532
rect 36988 45778 37044 45780
rect 36988 45726 36990 45778
rect 36990 45726 37042 45778
rect 37042 45726 37044 45778
rect 36988 45724 37044 45726
rect 36316 45612 36372 45668
rect 34860 45164 34916 45220
rect 34636 45106 34692 45108
rect 34636 45054 34638 45106
rect 34638 45054 34690 45106
rect 34690 45054 34692 45106
rect 34636 45052 34692 45054
rect 33964 44434 34020 44436
rect 33964 44382 33966 44434
rect 33966 44382 34018 44434
rect 34018 44382 34020 44434
rect 33964 44380 34020 44382
rect 34300 44882 34356 44884
rect 34300 44830 34302 44882
rect 34302 44830 34354 44882
rect 34354 44830 34356 44882
rect 34300 44828 34356 44830
rect 34188 44268 34244 44324
rect 33740 43762 33796 43764
rect 33740 43710 33742 43762
rect 33742 43710 33794 43762
rect 33794 43710 33796 43762
rect 33740 43708 33796 43710
rect 34188 43708 34244 43764
rect 35756 45106 35812 45108
rect 35756 45054 35758 45106
rect 35758 45054 35810 45106
rect 35810 45054 35812 45106
rect 35756 45052 35812 45054
rect 35420 44940 35476 44996
rect 35196 44714 35252 44716
rect 35196 44662 35198 44714
rect 35198 44662 35250 44714
rect 35250 44662 35252 44714
rect 35196 44660 35252 44662
rect 35300 44714 35356 44716
rect 35300 44662 35302 44714
rect 35302 44662 35354 44714
rect 35354 44662 35356 44714
rect 35300 44660 35356 44662
rect 35404 44714 35460 44716
rect 35404 44662 35406 44714
rect 35406 44662 35458 44714
rect 35458 44662 35460 44714
rect 35404 44660 35460 44662
rect 34860 44380 34916 44436
rect 35756 44322 35812 44324
rect 35756 44270 35758 44322
rect 35758 44270 35810 44322
rect 35810 44270 35812 44322
rect 35756 44268 35812 44270
rect 37660 49420 37716 49476
rect 37884 49420 37940 49476
rect 37548 48860 37604 48916
rect 38556 49756 38612 49812
rect 38220 49026 38276 49028
rect 38220 48974 38222 49026
rect 38222 48974 38274 49026
rect 38274 48974 38276 49026
rect 38220 48972 38276 48974
rect 37548 46396 37604 46452
rect 37324 45330 37380 45332
rect 37324 45278 37326 45330
rect 37326 45278 37378 45330
rect 37378 45278 37380 45330
rect 37324 45276 37380 45278
rect 37436 45106 37492 45108
rect 37436 45054 37438 45106
rect 37438 45054 37490 45106
rect 37490 45054 37492 45106
rect 37436 45052 37492 45054
rect 33180 42194 33236 42196
rect 33180 42142 33182 42194
rect 33182 42142 33234 42194
rect 33234 42142 33236 42194
rect 33180 42140 33236 42142
rect 33292 41746 33348 41748
rect 33292 41694 33294 41746
rect 33294 41694 33346 41746
rect 33346 41694 33348 41746
rect 33292 41692 33348 41694
rect 32172 41580 32228 41636
rect 32172 40236 32228 40292
rect 28028 37378 28084 37380
rect 28028 37326 28030 37378
rect 28030 37326 28082 37378
rect 28082 37326 28084 37378
rect 28028 37324 28084 37326
rect 28588 37938 28644 37940
rect 28588 37886 28590 37938
rect 28590 37886 28642 37938
rect 28642 37886 28644 37938
rect 28588 37884 28644 37886
rect 28476 37772 28532 37828
rect 28476 36204 28532 36260
rect 28140 36092 28196 36148
rect 28700 35196 28756 35252
rect 28364 34860 28420 34916
rect 28364 31948 28420 32004
rect 28364 31724 28420 31780
rect 28140 28812 28196 28868
rect 28252 31612 28308 31668
rect 28924 37266 28980 37268
rect 28924 37214 28926 37266
rect 28926 37214 28978 37266
rect 28978 37214 28980 37266
rect 28924 37212 28980 37214
rect 28924 29148 28980 29204
rect 28364 28812 28420 28868
rect 28252 28028 28308 28084
rect 28700 28476 28756 28532
rect 27468 27580 27524 27636
rect 27468 27132 27524 27188
rect 28588 27468 28644 27524
rect 28588 26962 28644 26964
rect 28588 26910 28590 26962
rect 28590 26910 28642 26962
rect 28642 26910 28644 26962
rect 28588 26908 28644 26910
rect 28700 27356 28756 27412
rect 28028 26178 28084 26180
rect 28028 26126 28030 26178
rect 28030 26126 28082 26178
rect 28082 26126 28084 26178
rect 28028 26124 28084 26126
rect 28812 26572 28868 26628
rect 29484 37884 29540 37940
rect 29260 37826 29316 37828
rect 29260 37774 29262 37826
rect 29262 37774 29314 37826
rect 29314 37774 29316 37826
rect 29260 37772 29316 37774
rect 29372 37490 29428 37492
rect 29372 37438 29374 37490
rect 29374 37438 29426 37490
rect 29426 37438 29428 37490
rect 29372 37436 29428 37438
rect 29148 36204 29204 36260
rect 30268 35308 30324 35364
rect 29148 34972 29204 35028
rect 29148 33068 29204 33124
rect 29260 35196 29316 35252
rect 29708 33346 29764 33348
rect 29708 33294 29710 33346
rect 29710 33294 29762 33346
rect 29762 33294 29764 33346
rect 29708 33292 29764 33294
rect 30380 34242 30436 34244
rect 30380 34190 30382 34242
rect 30382 34190 30434 34242
rect 30434 34190 30436 34242
rect 30380 34188 30436 34190
rect 30380 33852 30436 33908
rect 30268 33292 30324 33348
rect 32396 41298 32452 41300
rect 32396 41246 32398 41298
rect 32398 41246 32450 41298
rect 32450 41246 32452 41298
rect 32396 41244 32452 41246
rect 33516 41244 33572 41300
rect 33292 40236 33348 40292
rect 33964 43484 34020 43540
rect 34076 43372 34132 43428
rect 34860 43426 34916 43428
rect 34860 43374 34862 43426
rect 34862 43374 34914 43426
rect 34914 43374 34916 43426
rect 34860 43372 34916 43374
rect 35196 43146 35252 43148
rect 35196 43094 35198 43146
rect 35198 43094 35250 43146
rect 35250 43094 35252 43146
rect 35196 43092 35252 43094
rect 35300 43146 35356 43148
rect 35300 43094 35302 43146
rect 35302 43094 35354 43146
rect 35354 43094 35356 43146
rect 35300 43092 35356 43094
rect 35404 43146 35460 43148
rect 35404 43094 35406 43146
rect 35406 43094 35458 43146
rect 35458 43094 35460 43146
rect 35404 43092 35460 43094
rect 36428 42924 36484 42980
rect 36988 43260 37044 43316
rect 36988 42754 37044 42756
rect 36988 42702 36990 42754
rect 36990 42702 37042 42754
rect 37042 42702 37044 42754
rect 36988 42700 37044 42702
rect 38668 49084 38724 49140
rect 39788 49084 39844 49140
rect 38556 49026 38612 49028
rect 38556 48974 38558 49026
rect 38558 48974 38610 49026
rect 38610 48974 38612 49026
rect 38556 48972 38612 48974
rect 37996 48914 38052 48916
rect 37996 48862 37998 48914
rect 37998 48862 38050 48914
rect 38050 48862 38052 48914
rect 37996 48860 38052 48862
rect 38668 48860 38724 48916
rect 38444 48802 38500 48804
rect 38444 48750 38446 48802
rect 38446 48750 38498 48802
rect 38498 48750 38500 48802
rect 38444 48748 38500 48750
rect 37996 48188 38052 48244
rect 38556 47570 38612 47572
rect 38556 47518 38558 47570
rect 38558 47518 38610 47570
rect 38610 47518 38612 47570
rect 38556 47516 38612 47518
rect 38332 46562 38388 46564
rect 38332 46510 38334 46562
rect 38334 46510 38386 46562
rect 38386 46510 38388 46562
rect 38332 46508 38388 46510
rect 37884 45778 37940 45780
rect 37884 45726 37886 45778
rect 37886 45726 37938 45778
rect 37938 45726 37940 45778
rect 37884 45724 37940 45726
rect 38220 45890 38276 45892
rect 38220 45838 38222 45890
rect 38222 45838 38274 45890
rect 38274 45838 38276 45890
rect 38220 45836 38276 45838
rect 39004 48748 39060 48804
rect 38892 46674 38948 46676
rect 38892 46622 38894 46674
rect 38894 46622 38946 46674
rect 38946 46622 38948 46674
rect 38892 46620 38948 46622
rect 38780 46562 38836 46564
rect 38780 46510 38782 46562
rect 38782 46510 38834 46562
rect 38834 46510 38836 46562
rect 38780 46508 38836 46510
rect 38668 45724 38724 45780
rect 38780 45276 38836 45332
rect 38332 45218 38388 45220
rect 38332 45166 38334 45218
rect 38334 45166 38386 45218
rect 38386 45166 38388 45218
rect 38332 45164 38388 45166
rect 38444 45106 38500 45108
rect 38444 45054 38446 45106
rect 38446 45054 38498 45106
rect 38498 45054 38500 45106
rect 38444 45052 38500 45054
rect 38892 45218 38948 45220
rect 38892 45166 38894 45218
rect 38894 45166 38946 45218
rect 38946 45166 38948 45218
rect 38892 45164 38948 45166
rect 38668 44098 38724 44100
rect 38668 44046 38670 44098
rect 38670 44046 38722 44098
rect 38722 44046 38724 44098
rect 38668 44044 38724 44046
rect 40012 48972 40068 49028
rect 40348 48748 40404 48804
rect 40124 48076 40180 48132
rect 40012 47404 40068 47460
rect 40012 46620 40068 46676
rect 39564 45778 39620 45780
rect 39564 45726 39566 45778
rect 39566 45726 39618 45778
rect 39618 45726 39620 45778
rect 39564 45724 39620 45726
rect 39452 45218 39508 45220
rect 39452 45166 39454 45218
rect 39454 45166 39506 45218
rect 39506 45166 39508 45218
rect 39452 45164 39508 45166
rect 39564 44044 39620 44100
rect 38332 42924 38388 42980
rect 37772 42754 37828 42756
rect 37772 42702 37774 42754
rect 37774 42702 37826 42754
rect 37826 42702 37828 42754
rect 37772 42700 37828 42702
rect 34076 42476 34132 42532
rect 35196 41578 35252 41580
rect 35196 41526 35198 41578
rect 35198 41526 35250 41578
rect 35250 41526 35252 41578
rect 35196 41524 35252 41526
rect 35300 41578 35356 41580
rect 35300 41526 35302 41578
rect 35302 41526 35354 41578
rect 35354 41526 35356 41578
rect 35300 41524 35356 41526
rect 35404 41578 35460 41580
rect 35404 41526 35406 41578
rect 35406 41526 35458 41578
rect 35458 41526 35460 41578
rect 35404 41524 35460 41526
rect 35756 41244 35812 41300
rect 34300 41074 34356 41076
rect 34300 41022 34302 41074
rect 34302 41022 34354 41074
rect 34354 41022 34356 41074
rect 34300 41020 34356 41022
rect 35308 40514 35364 40516
rect 35308 40462 35310 40514
rect 35310 40462 35362 40514
rect 35362 40462 35364 40514
rect 35308 40460 35364 40462
rect 35196 40010 35252 40012
rect 35196 39958 35198 40010
rect 35198 39958 35250 40010
rect 35250 39958 35252 40010
rect 35196 39956 35252 39958
rect 35300 40010 35356 40012
rect 35300 39958 35302 40010
rect 35302 39958 35354 40010
rect 35354 39958 35356 40010
rect 35300 39956 35356 39958
rect 35404 40010 35460 40012
rect 35404 39958 35406 40010
rect 35406 39958 35458 40010
rect 35458 39958 35460 40010
rect 35404 39956 35460 39958
rect 36652 41244 36708 41300
rect 37100 41074 37156 41076
rect 37100 41022 37102 41074
rect 37102 41022 37154 41074
rect 37154 41022 37156 41074
rect 37100 41020 37156 41022
rect 36428 39564 36484 39620
rect 37100 39564 37156 39620
rect 36204 39228 36260 39284
rect 31948 37436 32004 37492
rect 34300 37938 34356 37940
rect 34300 37886 34302 37938
rect 34302 37886 34354 37938
rect 34354 37886 34356 37938
rect 34300 37884 34356 37886
rect 33740 37100 33796 37156
rect 29596 33122 29652 33124
rect 29596 33070 29598 33122
rect 29598 33070 29650 33122
rect 29650 33070 29652 33122
rect 29596 33068 29652 33070
rect 29260 32060 29316 32116
rect 30492 33122 30548 33124
rect 30492 33070 30494 33122
rect 30494 33070 30546 33122
rect 30546 33070 30548 33122
rect 30492 33068 30548 33070
rect 30380 32674 30436 32676
rect 30380 32622 30382 32674
rect 30382 32622 30434 32674
rect 30434 32622 30436 32674
rect 30380 32620 30436 32622
rect 30492 32562 30548 32564
rect 30492 32510 30494 32562
rect 30494 32510 30546 32562
rect 30546 32510 30548 32562
rect 30492 32508 30548 32510
rect 29932 31948 29988 32004
rect 30156 30492 30212 30548
rect 30940 33852 30996 33908
rect 32172 35026 32228 35028
rect 32172 34974 32174 35026
rect 32174 34974 32226 35026
rect 32226 34974 32228 35026
rect 32172 34972 32228 34974
rect 31276 33122 31332 33124
rect 31276 33070 31278 33122
rect 31278 33070 31330 33122
rect 31330 33070 31332 33122
rect 31276 33068 31332 33070
rect 30828 32562 30884 32564
rect 30828 32510 30830 32562
rect 30830 32510 30882 32562
rect 30882 32510 30884 32562
rect 30828 32508 30884 32510
rect 30940 32396 30996 32452
rect 31500 32620 31556 32676
rect 32284 32562 32340 32564
rect 32284 32510 32286 32562
rect 32286 32510 32338 32562
rect 32338 32510 32340 32562
rect 32284 32508 32340 32510
rect 30716 30492 30772 30548
rect 29372 30210 29428 30212
rect 29372 30158 29374 30210
rect 29374 30158 29426 30210
rect 29426 30158 29428 30210
rect 29372 30156 29428 30158
rect 29820 30156 29876 30212
rect 29036 28476 29092 28532
rect 29372 28866 29428 28868
rect 29372 28814 29374 28866
rect 29374 28814 29426 28866
rect 29426 28814 29428 28866
rect 29372 28812 29428 28814
rect 31164 30044 31220 30100
rect 30716 29986 30772 29988
rect 30716 29934 30718 29986
rect 30718 29934 30770 29986
rect 30770 29934 30772 29986
rect 30716 29932 30772 29934
rect 30380 28924 30436 28980
rect 30268 28476 30324 28532
rect 31164 29036 31220 29092
rect 29484 28418 29540 28420
rect 29484 28366 29486 28418
rect 29486 28366 29538 28418
rect 29538 28366 29540 28418
rect 29484 28364 29540 28366
rect 29708 27356 29764 27412
rect 29260 26962 29316 26964
rect 29260 26910 29262 26962
rect 29262 26910 29314 26962
rect 29314 26910 29316 26962
rect 29260 26908 29316 26910
rect 29372 26796 29428 26852
rect 29260 26572 29316 26628
rect 28924 26348 28980 26404
rect 30044 28364 30100 28420
rect 29932 26796 29988 26852
rect 30604 28476 30660 28532
rect 31052 28476 31108 28532
rect 30380 28364 30436 28420
rect 30940 28418 30996 28420
rect 30940 28366 30942 28418
rect 30942 28366 30994 28418
rect 30994 28366 30996 28418
rect 30940 28364 30996 28366
rect 30604 27186 30660 27188
rect 30604 27134 30606 27186
rect 30606 27134 30658 27186
rect 30658 27134 30660 27186
rect 30604 27132 30660 27134
rect 31500 29932 31556 29988
rect 30940 27020 30996 27076
rect 30268 26962 30324 26964
rect 30268 26910 30270 26962
rect 30270 26910 30322 26962
rect 30322 26910 30324 26962
rect 30268 26908 30324 26910
rect 29708 26684 29764 26740
rect 30268 26684 30324 26740
rect 29484 26178 29540 26180
rect 29484 26126 29486 26178
rect 29486 26126 29538 26178
rect 29538 26126 29540 26178
rect 29484 26124 29540 26126
rect 30268 26124 30324 26180
rect 30828 26402 30884 26404
rect 30828 26350 30830 26402
rect 30830 26350 30882 26402
rect 30882 26350 30884 26402
rect 30828 26348 30884 26350
rect 31164 26572 31220 26628
rect 31500 26684 31556 26740
rect 31500 26402 31556 26404
rect 31500 26350 31502 26402
rect 31502 26350 31554 26402
rect 31554 26350 31556 26402
rect 31500 26348 31556 26350
rect 30044 25452 30100 25508
rect 29820 25394 29876 25396
rect 29820 25342 29822 25394
rect 29822 25342 29874 25394
rect 29874 25342 29876 25394
rect 29820 25340 29876 25342
rect 29708 25116 29764 25172
rect 26796 24946 26852 24948
rect 26796 24894 26798 24946
rect 26798 24894 26850 24946
rect 26850 24894 26852 24946
rect 26796 24892 26852 24894
rect 26460 22204 26516 22260
rect 25452 17500 25508 17556
rect 26348 21868 26404 21924
rect 25900 17612 25956 17668
rect 24108 15036 24164 15092
rect 25564 16716 25620 16772
rect 25900 16604 25956 16660
rect 25340 15260 25396 15316
rect 26684 23436 26740 23492
rect 29036 25004 29092 25060
rect 28028 23324 28084 23380
rect 26908 22876 26964 22932
rect 26684 22428 26740 22484
rect 26572 22092 26628 22148
rect 26908 21980 26964 22036
rect 23996 12850 24052 12852
rect 23996 12798 23998 12850
rect 23998 12798 24050 12850
rect 24050 12798 24052 12850
rect 23996 12796 24052 12798
rect 23884 12178 23940 12180
rect 23884 12126 23886 12178
rect 23886 12126 23938 12178
rect 23938 12126 23940 12178
rect 23884 12124 23940 12126
rect 24220 12178 24276 12180
rect 24220 12126 24222 12178
rect 24222 12126 24274 12178
rect 24274 12126 24276 12178
rect 24220 12124 24276 12126
rect 25340 13634 25396 13636
rect 25340 13582 25342 13634
rect 25342 13582 25394 13634
rect 25394 13582 25396 13634
rect 25340 13580 25396 13582
rect 25228 13356 25284 13412
rect 25228 12348 25284 12404
rect 25116 12124 25172 12180
rect 24780 11170 24836 11172
rect 24780 11118 24782 11170
rect 24782 11118 24834 11170
rect 24834 11118 24836 11170
rect 24780 11116 24836 11118
rect 20972 8428 21028 8484
rect 20524 8258 20580 8260
rect 20524 8206 20526 8258
rect 20526 8206 20578 8258
rect 20578 8206 20580 8258
rect 20524 8204 20580 8206
rect 20412 8146 20468 8148
rect 20412 8094 20414 8146
rect 20414 8094 20466 8146
rect 20466 8094 20468 8146
rect 20412 8092 20468 8094
rect 19628 7586 19684 7588
rect 19628 7534 19630 7586
rect 19630 7534 19682 7586
rect 19682 7534 19684 7586
rect 19628 7532 19684 7534
rect 20748 7980 20804 8036
rect 20300 7868 20356 7924
rect 19516 7420 19572 7476
rect 19852 7474 19908 7476
rect 19852 7422 19854 7474
rect 19854 7422 19906 7474
rect 19906 7422 19908 7474
rect 19852 7420 19908 7422
rect 19516 6076 19572 6132
rect 19964 7362 20020 7364
rect 19964 7310 19966 7362
rect 19966 7310 20018 7362
rect 20018 7310 20020 7362
rect 19964 7308 20020 7310
rect 17388 5852 17444 5908
rect 15260 5628 15316 5684
rect 18844 5682 18900 5684
rect 18844 5630 18846 5682
rect 18846 5630 18898 5682
rect 18898 5630 18900 5682
rect 18844 5628 18900 5630
rect 14700 5068 14756 5124
rect 16828 5068 16884 5124
rect 17836 5122 17892 5124
rect 17836 5070 17838 5122
rect 17838 5070 17890 5122
rect 17890 5070 17892 5122
rect 17836 5068 17892 5070
rect 14364 4396 14420 4452
rect 14924 4450 14980 4452
rect 14924 4398 14926 4450
rect 14926 4398 14978 4450
rect 14978 4398 14980 4450
rect 14924 4396 14980 4398
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19740 6130 19796 6132
rect 19740 6078 19742 6130
rect 19742 6078 19794 6130
rect 19794 6078 19796 6130
rect 19740 6076 19796 6078
rect 20860 7698 20916 7700
rect 20860 7646 20862 7698
rect 20862 7646 20914 7698
rect 20914 7646 20916 7698
rect 20860 7644 20916 7646
rect 20300 7420 20356 7476
rect 20636 7362 20692 7364
rect 20636 7310 20638 7362
rect 20638 7310 20690 7362
rect 20690 7310 20692 7362
rect 20636 7308 20692 7310
rect 20748 6748 20804 6804
rect 20188 6076 20244 6132
rect 19964 6018 20020 6020
rect 19964 5966 19966 6018
rect 19966 5966 20018 6018
rect 20018 5966 20020 6018
rect 19964 5964 20020 5966
rect 19628 5906 19684 5908
rect 19628 5854 19630 5906
rect 19630 5854 19682 5906
rect 19682 5854 19684 5906
rect 19628 5852 19684 5854
rect 20300 5964 20356 6020
rect 19180 5346 19236 5348
rect 19180 5294 19182 5346
rect 19182 5294 19234 5346
rect 19234 5294 19236 5346
rect 19180 5292 19236 5294
rect 18956 5068 19012 5124
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 21980 8204 22036 8260
rect 22204 8876 22260 8932
rect 22652 8258 22708 8260
rect 22652 8206 22654 8258
rect 22654 8206 22706 8258
rect 22706 8206 22708 8258
rect 22652 8204 22708 8206
rect 22092 8034 22148 8036
rect 22092 7982 22094 8034
rect 22094 7982 22146 8034
rect 22146 7982 22148 8034
rect 22092 7980 22148 7982
rect 21644 6412 21700 6468
rect 23100 7980 23156 8036
rect 22428 7868 22484 7924
rect 23548 7698 23604 7700
rect 23548 7646 23550 7698
rect 23550 7646 23602 7698
rect 23602 7646 23604 7698
rect 23548 7644 23604 7646
rect 22316 7474 22372 7476
rect 22316 7422 22318 7474
rect 22318 7422 22370 7474
rect 22370 7422 22372 7474
rect 22316 7420 22372 7422
rect 25564 12348 25620 12404
rect 25340 11116 25396 11172
rect 25116 9884 25172 9940
rect 26124 14306 26180 14308
rect 26124 14254 26126 14306
rect 26126 14254 26178 14306
rect 26178 14254 26180 14306
rect 26124 14252 26180 14254
rect 26572 14306 26628 14308
rect 26572 14254 26574 14306
rect 26574 14254 26626 14306
rect 26626 14254 26628 14306
rect 26572 14252 26628 14254
rect 26460 13580 26516 13636
rect 26348 13356 26404 13412
rect 27020 21644 27076 21700
rect 28252 22370 28308 22372
rect 28252 22318 28254 22370
rect 28254 22318 28306 22370
rect 28306 22318 28308 22370
rect 28252 22316 28308 22318
rect 27692 21644 27748 21700
rect 27020 20802 27076 20804
rect 27020 20750 27022 20802
rect 27022 20750 27074 20802
rect 27074 20750 27076 20802
rect 27020 20748 27076 20750
rect 27916 20802 27972 20804
rect 27916 20750 27918 20802
rect 27918 20750 27970 20802
rect 27970 20750 27972 20802
rect 27916 20748 27972 20750
rect 27692 20636 27748 20692
rect 27244 20076 27300 20132
rect 27916 20412 27972 20468
rect 28476 20802 28532 20804
rect 28476 20750 28478 20802
rect 28478 20750 28530 20802
rect 28530 20750 28532 20802
rect 28476 20748 28532 20750
rect 28364 20412 28420 20468
rect 28028 20018 28084 20020
rect 28028 19966 28030 20018
rect 28030 19966 28082 20018
rect 28082 19966 28084 20018
rect 28028 19964 28084 19966
rect 28476 20076 28532 20132
rect 28140 19852 28196 19908
rect 27916 14252 27972 14308
rect 27692 13692 27748 13748
rect 26796 13634 26852 13636
rect 26796 13582 26798 13634
rect 26798 13582 26850 13634
rect 26850 13582 26852 13634
rect 26796 13580 26852 13582
rect 26684 13020 26740 13076
rect 27692 13020 27748 13076
rect 27132 12348 27188 12404
rect 25788 9884 25844 9940
rect 25564 8204 25620 8260
rect 24780 7980 24836 8036
rect 25900 8204 25956 8260
rect 25676 7532 25732 7588
rect 26236 11282 26292 11284
rect 26236 11230 26238 11282
rect 26238 11230 26290 11282
rect 26290 11230 26292 11282
rect 26236 11228 26292 11230
rect 26684 11228 26740 11284
rect 26460 9938 26516 9940
rect 26460 9886 26462 9938
rect 26462 9886 26514 9938
rect 26514 9886 26516 9938
rect 26460 9884 26516 9886
rect 26572 8428 26628 8484
rect 26348 8034 26404 8036
rect 26348 7982 26350 8034
rect 26350 7982 26402 8034
rect 26402 7982 26404 8034
rect 26348 7980 26404 7982
rect 23548 7084 23604 7140
rect 22876 6412 22932 6468
rect 22428 6188 22484 6244
rect 21756 6130 21812 6132
rect 21756 6078 21758 6130
rect 21758 6078 21810 6130
rect 21810 6078 21812 6130
rect 21756 6076 21812 6078
rect 21308 5964 21364 6020
rect 21420 5906 21476 5908
rect 21420 5854 21422 5906
rect 21422 5854 21474 5906
rect 21474 5854 21476 5906
rect 21420 5852 21476 5854
rect 24444 6412 24500 6468
rect 22652 5906 22708 5908
rect 22652 5854 22654 5906
rect 22654 5854 22706 5906
rect 22706 5854 22708 5906
rect 22652 5852 22708 5854
rect 21532 5292 21588 5348
rect 22540 5068 22596 5124
rect 21644 4338 21700 4340
rect 21644 4286 21646 4338
rect 21646 4286 21698 4338
rect 21698 4286 21700 4338
rect 21644 4284 21700 4286
rect 25788 7084 25844 7140
rect 25228 5068 25284 5124
rect 25788 5122 25844 5124
rect 25788 5070 25790 5122
rect 25790 5070 25842 5122
rect 25842 5070 25844 5122
rect 25788 5068 25844 5070
rect 26124 5122 26180 5124
rect 26124 5070 26126 5122
rect 26126 5070 26178 5122
rect 26178 5070 26180 5122
rect 26124 5068 26180 5070
rect 24668 4284 24724 4340
rect 25228 4338 25284 4340
rect 25228 4286 25230 4338
rect 25230 4286 25282 4338
rect 25282 4286 25284 4338
rect 25228 4284 25284 4286
rect 10780 3500 10836 3556
rect 7196 3388 7252 3444
rect 10108 3442 10164 3444
rect 10108 3390 10110 3442
rect 10110 3390 10162 3442
rect 10162 3390 10164 3442
rect 10108 3388 10164 3390
rect 11900 3612 11956 3668
rect 12460 3666 12516 3668
rect 12460 3614 12462 3666
rect 12462 3614 12514 3666
rect 12514 3614 12516 3666
rect 12460 3612 12516 3614
rect 28812 24722 28868 24724
rect 28812 24670 28814 24722
rect 28814 24670 28866 24722
rect 28866 24670 28868 24722
rect 28812 24668 28868 24670
rect 29148 24946 29204 24948
rect 29148 24894 29150 24946
rect 29150 24894 29202 24946
rect 29202 24894 29204 24946
rect 29148 24892 29204 24894
rect 29372 23042 29428 23044
rect 29372 22990 29374 23042
rect 29374 22990 29426 23042
rect 29426 22990 29428 23042
rect 29372 22988 29428 22990
rect 29148 22370 29204 22372
rect 29148 22318 29150 22370
rect 29150 22318 29202 22370
rect 29202 22318 29204 22370
rect 29148 22316 29204 22318
rect 29484 22258 29540 22260
rect 29484 22206 29486 22258
rect 29486 22206 29538 22258
rect 29538 22206 29540 22258
rect 29484 22204 29540 22206
rect 30380 25282 30436 25284
rect 30380 25230 30382 25282
rect 30382 25230 30434 25282
rect 30434 25230 30436 25282
rect 30380 25228 30436 25230
rect 31164 25394 31220 25396
rect 31164 25342 31166 25394
rect 31166 25342 31218 25394
rect 31218 25342 31220 25394
rect 31164 25340 31220 25342
rect 30380 22988 30436 23044
rect 29036 20690 29092 20692
rect 29036 20638 29038 20690
rect 29038 20638 29090 20690
rect 29090 20638 29092 20690
rect 29036 20636 29092 20638
rect 30268 20802 30324 20804
rect 30268 20750 30270 20802
rect 30270 20750 30322 20802
rect 30322 20750 30324 20802
rect 30268 20748 30324 20750
rect 28812 20018 28868 20020
rect 28812 19966 28814 20018
rect 28814 19966 28866 20018
rect 28866 19966 28868 20018
rect 28812 19964 28868 19966
rect 28700 19628 28756 19684
rect 29260 19628 29316 19684
rect 30044 20242 30100 20244
rect 30044 20190 30046 20242
rect 30046 20190 30098 20242
rect 30098 20190 30100 20242
rect 30044 20188 30100 20190
rect 29596 17666 29652 17668
rect 29596 17614 29598 17666
rect 29598 17614 29650 17666
rect 29650 17614 29652 17666
rect 29596 17612 29652 17614
rect 30604 21644 30660 21700
rect 30940 23714 30996 23716
rect 30940 23662 30942 23714
rect 30942 23662 30994 23714
rect 30994 23662 30996 23714
rect 30940 23660 30996 23662
rect 30828 22204 30884 22260
rect 30828 21868 30884 21924
rect 30940 21644 30996 21700
rect 30828 21532 30884 21588
rect 30492 20188 30548 20244
rect 31388 24780 31444 24836
rect 31164 24722 31220 24724
rect 31164 24670 31166 24722
rect 31166 24670 31218 24722
rect 31218 24670 31220 24722
rect 31164 24668 31220 24670
rect 31276 24444 31332 24500
rect 31948 32450 32004 32452
rect 31948 32398 31950 32450
rect 31950 32398 32002 32450
rect 32002 32398 32004 32450
rect 31948 32396 32004 32398
rect 31948 31554 32004 31556
rect 31948 31502 31950 31554
rect 31950 31502 32002 31554
rect 32002 31502 32004 31554
rect 31948 31500 32004 31502
rect 31836 30098 31892 30100
rect 31836 30046 31838 30098
rect 31838 30046 31890 30098
rect 31890 30046 31892 30098
rect 31836 30044 31892 30046
rect 31836 27970 31892 27972
rect 31836 27918 31838 27970
rect 31838 27918 31890 27970
rect 31890 27918 31892 27970
rect 31836 27916 31892 27918
rect 31836 27186 31892 27188
rect 31836 27134 31838 27186
rect 31838 27134 31890 27186
rect 31890 27134 31892 27186
rect 31836 27132 31892 27134
rect 31724 26796 31780 26852
rect 31836 25340 31892 25396
rect 31052 19628 31108 19684
rect 30716 18956 30772 19012
rect 30044 17666 30100 17668
rect 30044 17614 30046 17666
rect 30046 17614 30098 17666
rect 30098 17614 30100 17666
rect 30044 17612 30100 17614
rect 29820 16156 29876 16212
rect 30940 18844 30996 18900
rect 31164 19404 31220 19460
rect 31052 18172 31108 18228
rect 31164 19068 31220 19124
rect 29260 15148 29316 15204
rect 30940 15036 30996 15092
rect 31500 23378 31556 23380
rect 31500 23326 31502 23378
rect 31502 23326 31554 23378
rect 31554 23326 31556 23378
rect 31500 23324 31556 23326
rect 31612 21532 31668 21588
rect 31724 21420 31780 21476
rect 31612 19852 31668 19908
rect 32732 35308 32788 35364
rect 33068 35308 33124 35364
rect 33516 35308 33572 35364
rect 33068 33852 33124 33908
rect 33180 34300 33236 34356
rect 33852 34300 33908 34356
rect 33180 33292 33236 33348
rect 32844 33122 32900 33124
rect 32844 33070 32846 33122
rect 32846 33070 32898 33122
rect 32898 33070 32900 33122
rect 32844 33068 32900 33070
rect 32508 31724 32564 31780
rect 33180 32508 33236 32564
rect 32396 31500 32452 31556
rect 33852 33346 33908 33348
rect 33852 33294 33854 33346
rect 33854 33294 33906 33346
rect 33906 33294 33908 33346
rect 33852 33292 33908 33294
rect 33740 33234 33796 33236
rect 33740 33182 33742 33234
rect 33742 33182 33794 33234
rect 33794 33182 33796 33234
rect 33740 33180 33796 33182
rect 34300 33234 34356 33236
rect 34300 33182 34302 33234
rect 34302 33182 34354 33234
rect 34354 33182 34356 33234
rect 34300 33180 34356 33182
rect 33516 32508 33572 32564
rect 33740 32060 33796 32116
rect 33516 31836 33572 31892
rect 33292 31500 33348 31556
rect 32396 30156 32452 30212
rect 32396 29372 32452 29428
rect 33516 31500 33572 31556
rect 33292 30268 33348 30324
rect 32172 28812 32228 28868
rect 32284 25116 32340 25172
rect 34412 32450 34468 32452
rect 34412 32398 34414 32450
rect 34414 32398 34466 32450
rect 34466 32398 34468 32450
rect 34412 32396 34468 32398
rect 34300 32060 34356 32116
rect 34748 31836 34804 31892
rect 34636 31500 34692 31556
rect 33852 31276 33908 31332
rect 34748 31276 34804 31332
rect 33740 30828 33796 30884
rect 33628 29986 33684 29988
rect 33628 29934 33630 29986
rect 33630 29934 33682 29986
rect 33682 29934 33684 29986
rect 33628 29932 33684 29934
rect 34636 30210 34692 30212
rect 34636 30158 34638 30210
rect 34638 30158 34690 30210
rect 34690 30158 34692 30210
rect 34636 30156 34692 30158
rect 33964 29986 34020 29988
rect 33964 29934 33966 29986
rect 33966 29934 34018 29986
rect 34018 29934 34020 29986
rect 33964 29932 34020 29934
rect 33740 29596 33796 29652
rect 34412 29932 34468 29988
rect 34188 28476 34244 28532
rect 34076 28364 34132 28420
rect 34748 28364 34804 28420
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 37212 39228 37268 39284
rect 36428 37154 36484 37156
rect 36428 37102 36430 37154
rect 36430 37102 36482 37154
rect 36482 37102 36484 37154
rect 36428 37100 36484 37102
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 36204 36370 36260 36372
rect 36204 36318 36206 36370
rect 36206 36318 36258 36370
rect 36258 36318 36260 36370
rect 36204 36316 36260 36318
rect 35756 35868 35812 35924
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35756 34972 35812 35028
rect 38668 42978 38724 42980
rect 38668 42926 38670 42978
rect 38670 42926 38722 42978
rect 38722 42926 38724 42978
rect 38668 42924 38724 42926
rect 38780 42700 38836 42756
rect 39004 42642 39060 42644
rect 39004 42590 39006 42642
rect 39006 42590 39058 42642
rect 39058 42590 39060 42642
rect 39004 42588 39060 42590
rect 38444 42194 38500 42196
rect 38444 42142 38446 42194
rect 38446 42142 38498 42194
rect 38498 42142 38500 42194
rect 38444 42140 38500 42142
rect 38892 40626 38948 40628
rect 38892 40574 38894 40626
rect 38894 40574 38946 40626
rect 38946 40574 38948 40626
rect 38892 40572 38948 40574
rect 38108 40460 38164 40516
rect 38332 40236 38388 40292
rect 37548 38050 37604 38052
rect 37548 37998 37550 38050
rect 37550 37998 37602 38050
rect 37602 37998 37604 38050
rect 37548 37996 37604 37998
rect 37100 37938 37156 37940
rect 37100 37886 37102 37938
rect 37102 37886 37154 37938
rect 37154 37886 37156 37938
rect 37100 37884 37156 37886
rect 37100 37154 37156 37156
rect 37100 37102 37102 37154
rect 37102 37102 37154 37154
rect 37154 37102 37156 37154
rect 37100 37100 37156 37102
rect 37548 37100 37604 37156
rect 38220 36540 38276 36596
rect 37324 36316 37380 36372
rect 36540 34972 36596 35028
rect 36204 34914 36260 34916
rect 36204 34862 36206 34914
rect 36206 34862 36258 34914
rect 36258 34862 36260 34914
rect 36204 34860 36260 34862
rect 35980 34636 36036 34692
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 37100 34690 37156 34692
rect 37100 34638 37102 34690
rect 37102 34638 37154 34690
rect 37154 34638 37156 34690
rect 37100 34636 37156 34638
rect 38444 39730 38500 39732
rect 38444 39678 38446 39730
rect 38446 39678 38498 39730
rect 38498 39678 38500 39730
rect 38444 39676 38500 39678
rect 38556 39228 38612 39284
rect 38780 37100 38836 37156
rect 39004 36652 39060 36708
rect 38892 36594 38948 36596
rect 38892 36542 38894 36594
rect 38894 36542 38946 36594
rect 38946 36542 38948 36594
rect 38892 36540 38948 36542
rect 39340 42700 39396 42756
rect 39228 39340 39284 39396
rect 38220 35698 38276 35700
rect 38220 35646 38222 35698
rect 38222 35646 38274 35698
rect 38274 35646 38276 35698
rect 38220 35644 38276 35646
rect 36988 34412 37044 34468
rect 35756 33180 35812 33236
rect 35868 33852 35924 33908
rect 35308 32562 35364 32564
rect 35308 32510 35310 32562
rect 35310 32510 35362 32562
rect 35362 32510 35364 32562
rect 35308 32508 35364 32510
rect 35532 32284 35588 32340
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35084 31836 35140 31892
rect 34860 27916 34916 27972
rect 34972 30828 35028 30884
rect 34748 27858 34804 27860
rect 34748 27806 34750 27858
rect 34750 27806 34802 27858
rect 34802 27806 34804 27858
rect 34748 27804 34804 27806
rect 33740 27020 33796 27076
rect 33516 26236 33572 26292
rect 32284 24834 32340 24836
rect 32284 24782 32286 24834
rect 32286 24782 32338 24834
rect 32338 24782 32340 24834
rect 32284 24780 32340 24782
rect 32172 24668 32228 24724
rect 32172 24498 32228 24500
rect 32172 24446 32174 24498
rect 32174 24446 32226 24498
rect 32226 24446 32228 24498
rect 32172 24444 32228 24446
rect 33292 24498 33348 24500
rect 33292 24446 33294 24498
rect 33294 24446 33346 24498
rect 33346 24446 33348 24498
rect 33292 24444 33348 24446
rect 33516 24892 33572 24948
rect 33628 25564 33684 25620
rect 33404 23996 33460 24052
rect 32060 20748 32116 20804
rect 31612 19180 31668 19236
rect 33628 23548 33684 23604
rect 33180 21644 33236 21700
rect 33404 21474 33460 21476
rect 33404 21422 33406 21474
rect 33406 21422 33458 21474
rect 33458 21422 33460 21474
rect 33404 21420 33460 21422
rect 33964 26684 34020 26740
rect 34748 27468 34804 27524
rect 34076 26908 34132 26964
rect 33852 26572 33908 26628
rect 33852 24722 33908 24724
rect 33852 24670 33854 24722
rect 33854 24670 33906 24722
rect 33906 24670 33908 24722
rect 33852 24668 33908 24670
rect 34748 26572 34804 26628
rect 35196 31554 35252 31556
rect 35196 31502 35198 31554
rect 35198 31502 35250 31554
rect 35250 31502 35252 31554
rect 35196 31500 35252 31502
rect 35196 30882 35252 30884
rect 35196 30830 35198 30882
rect 35198 30830 35250 30882
rect 35250 30830 35252 30882
rect 35196 30828 35252 30830
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35980 32450 36036 32452
rect 35980 32398 35982 32450
rect 35982 32398 36034 32450
rect 36034 32398 36036 32450
rect 35980 32396 36036 32398
rect 38332 34914 38388 34916
rect 38332 34862 38334 34914
rect 38334 34862 38386 34914
rect 38386 34862 38388 34914
rect 38332 34860 38388 34862
rect 37884 34412 37940 34468
rect 37100 31778 37156 31780
rect 37100 31726 37102 31778
rect 37102 31726 37154 31778
rect 37154 31726 37156 31778
rect 37100 31724 37156 31726
rect 37100 31276 37156 31332
rect 36988 31164 37044 31220
rect 36204 30828 36260 30884
rect 35084 29932 35140 29988
rect 35532 30380 35588 30436
rect 35532 30210 35588 30212
rect 35532 30158 35534 30210
rect 35534 30158 35586 30210
rect 35586 30158 35588 30210
rect 35532 30156 35588 30158
rect 38892 35922 38948 35924
rect 38892 35870 38894 35922
rect 38894 35870 38946 35922
rect 38946 35870 38948 35922
rect 38892 35868 38948 35870
rect 38892 34130 38948 34132
rect 38892 34078 38894 34130
rect 38894 34078 38946 34130
rect 38946 34078 38948 34130
rect 38892 34076 38948 34078
rect 39340 36204 39396 36260
rect 39340 35980 39396 36036
rect 39340 34972 39396 35028
rect 39452 33292 39508 33348
rect 38780 32562 38836 32564
rect 38780 32510 38782 32562
rect 38782 32510 38834 32562
rect 38834 32510 38836 32562
rect 38780 32508 38836 32510
rect 37436 32172 37492 32228
rect 36540 30882 36596 30884
rect 36540 30830 36542 30882
rect 36542 30830 36594 30882
rect 36594 30830 36596 30882
rect 36540 30828 36596 30830
rect 35756 29820 35812 29876
rect 36428 29820 36484 29876
rect 36316 29372 36372 29428
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27804 35252 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 35308 27186 35364 27188
rect 35308 27134 35310 27186
rect 35310 27134 35362 27186
rect 35362 27134 35364 27186
rect 35308 27132 35364 27134
rect 35196 26572 35252 26628
rect 35308 26684 35364 26740
rect 34188 24444 34244 24500
rect 34636 23548 34692 23604
rect 36204 28700 36260 28756
rect 36092 27858 36148 27860
rect 36092 27806 36094 27858
rect 36094 27806 36146 27858
rect 36146 27806 36148 27858
rect 36092 27804 36148 27806
rect 36428 28476 36484 28532
rect 36428 28082 36484 28084
rect 36428 28030 36430 28082
rect 36430 28030 36482 28082
rect 36482 28030 36484 28082
rect 36428 28028 36484 28030
rect 36988 29708 37044 29764
rect 36316 27692 36372 27748
rect 35756 27074 35812 27076
rect 35756 27022 35758 27074
rect 35758 27022 35810 27074
rect 35810 27022 35812 27074
rect 35756 27020 35812 27022
rect 36092 26908 36148 26964
rect 35756 26572 35812 26628
rect 35980 26684 36036 26740
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 35420 25506 35476 25508
rect 35420 25454 35422 25506
rect 35422 25454 35474 25506
rect 35474 25454 35476 25506
rect 35420 25452 35476 25454
rect 34860 24444 34916 24500
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 35196 24108 35252 24164
rect 34972 23660 35028 23716
rect 33964 22370 34020 22372
rect 33964 22318 33966 22370
rect 33966 22318 34018 22370
rect 34018 22318 34020 22370
rect 33964 22316 34020 22318
rect 33964 21868 34020 21924
rect 34860 22092 34916 22148
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 35420 22258 35476 22260
rect 35420 22206 35422 22258
rect 35422 22206 35474 22258
rect 35474 22206 35476 22258
rect 35420 22204 35476 22206
rect 36204 25564 36260 25620
rect 36316 25452 36372 25508
rect 36652 28588 36708 28644
rect 36652 27132 36708 27188
rect 36764 27858 36820 27860
rect 36764 27806 36766 27858
rect 36766 27806 36818 27858
rect 36818 27806 36820 27858
rect 36764 27804 36820 27806
rect 36540 26796 36596 26852
rect 36652 24444 36708 24500
rect 36428 22988 36484 23044
rect 36652 23154 36708 23156
rect 36652 23102 36654 23154
rect 36654 23102 36706 23154
rect 36706 23102 36708 23154
rect 36652 23100 36708 23102
rect 35308 22146 35364 22148
rect 35308 22094 35310 22146
rect 35310 22094 35362 22146
rect 35362 22094 35364 22146
rect 35308 22092 35364 22094
rect 35308 21756 35364 21812
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 32508 19292 32564 19348
rect 32172 19234 32228 19236
rect 32172 19182 32174 19234
rect 32174 19182 32226 19234
rect 32226 19182 32228 19234
rect 32172 19180 32228 19182
rect 33292 19234 33348 19236
rect 33292 19182 33294 19234
rect 33294 19182 33346 19234
rect 33346 19182 33348 19234
rect 33292 19180 33348 19182
rect 31836 19122 31892 19124
rect 31836 19070 31838 19122
rect 31838 19070 31890 19122
rect 31890 19070 31892 19122
rect 31836 19068 31892 19070
rect 32844 19122 32900 19124
rect 32844 19070 32846 19122
rect 32846 19070 32898 19122
rect 32898 19070 32900 19122
rect 32844 19068 32900 19070
rect 32620 19010 32676 19012
rect 32620 18958 32622 19010
rect 32622 18958 32674 19010
rect 32674 18958 32676 19010
rect 32620 18956 32676 18958
rect 31276 18844 31332 18900
rect 32732 17388 32788 17444
rect 33964 19010 34020 19012
rect 33964 18958 33966 19010
rect 33966 18958 34018 19010
rect 34018 18958 34020 19010
rect 33964 18956 34020 18958
rect 32956 17500 33012 17556
rect 33404 17554 33460 17556
rect 33404 17502 33406 17554
rect 33406 17502 33458 17554
rect 33458 17502 33460 17554
rect 33404 17500 33460 17502
rect 33516 17442 33572 17444
rect 33516 17390 33518 17442
rect 33518 17390 33570 17442
rect 33570 17390 33572 17442
rect 33516 17388 33572 17390
rect 32956 17052 33012 17108
rect 32844 16940 32900 16996
rect 31388 15538 31444 15540
rect 31388 15486 31390 15538
rect 31390 15486 31442 15538
rect 31442 15486 31444 15538
rect 31388 15484 31444 15486
rect 32396 15538 32452 15540
rect 32396 15486 32398 15538
rect 32398 15486 32450 15538
rect 32450 15486 32452 15538
rect 32396 15484 32452 15486
rect 31612 15036 31668 15092
rect 31276 14418 31332 14420
rect 31276 14366 31278 14418
rect 31278 14366 31330 14418
rect 31330 14366 31332 14418
rect 31276 14364 31332 14366
rect 31388 14306 31444 14308
rect 31388 14254 31390 14306
rect 31390 14254 31442 14306
rect 31442 14254 31444 14306
rect 31388 14252 31444 14254
rect 31164 13804 31220 13860
rect 32172 15036 32228 15092
rect 31836 13858 31892 13860
rect 31836 13806 31838 13858
rect 31838 13806 31890 13858
rect 31890 13806 31892 13858
rect 31836 13804 31892 13806
rect 32508 14700 32564 14756
rect 32284 14418 32340 14420
rect 32284 14366 32286 14418
rect 32286 14366 32338 14418
rect 32338 14366 32340 14418
rect 32284 14364 32340 14366
rect 32172 14252 32228 14308
rect 32396 14140 32452 14196
rect 31948 13692 32004 13748
rect 32508 13916 32564 13972
rect 31052 13244 31108 13300
rect 33404 16940 33460 16996
rect 34300 19292 34356 19348
rect 34636 19122 34692 19124
rect 34636 19070 34638 19122
rect 34638 19070 34690 19122
rect 34690 19070 34692 19122
rect 34636 19068 34692 19070
rect 34412 19010 34468 19012
rect 34412 18958 34414 19010
rect 34414 18958 34466 19010
rect 34466 18958 34468 19010
rect 34412 18956 34468 18958
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 34860 19292 34916 19348
rect 35308 19180 35364 19236
rect 35196 19122 35252 19124
rect 35196 19070 35198 19122
rect 35198 19070 35250 19122
rect 35250 19070 35252 19122
rect 35196 19068 35252 19070
rect 34972 18396 35028 18452
rect 34748 17500 34804 17556
rect 36428 18508 36484 18564
rect 36092 18450 36148 18452
rect 36092 18398 36094 18450
rect 36094 18398 36146 18450
rect 36146 18398 36148 18450
rect 36092 18396 36148 18398
rect 35420 18284 35476 18340
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 35084 17388 35140 17444
rect 36316 17442 36372 17444
rect 36316 17390 36318 17442
rect 36318 17390 36370 17442
rect 36370 17390 36372 17442
rect 36316 17388 36372 17390
rect 34188 16940 34244 16996
rect 33516 16828 33572 16884
rect 34300 16882 34356 16884
rect 34300 16830 34302 16882
rect 34302 16830 34354 16882
rect 34354 16830 34356 16882
rect 34300 16828 34356 16830
rect 33964 15202 34020 15204
rect 33964 15150 33966 15202
rect 33966 15150 34018 15202
rect 34018 15150 34020 15202
rect 33964 15148 34020 15150
rect 33068 14754 33124 14756
rect 33068 14702 33070 14754
rect 33070 14702 33122 14754
rect 33122 14702 33124 14754
rect 33068 14700 33124 14702
rect 33628 14700 33684 14756
rect 33180 14418 33236 14420
rect 33180 14366 33182 14418
rect 33182 14366 33234 14418
rect 33234 14366 33236 14418
rect 33180 14364 33236 14366
rect 33068 14306 33124 14308
rect 33068 14254 33070 14306
rect 33070 14254 33122 14306
rect 33122 14254 33124 14306
rect 33068 14252 33124 14254
rect 32956 13916 33012 13972
rect 33180 13804 33236 13860
rect 35308 17052 35364 17108
rect 35420 16994 35476 16996
rect 35420 16942 35422 16994
rect 35422 16942 35474 16994
rect 35474 16942 35476 16994
rect 35420 16940 35476 16942
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 34748 16268 34804 16324
rect 36316 16044 36372 16100
rect 36428 16716 36484 16772
rect 34524 15260 34580 15316
rect 34860 15986 34916 15988
rect 34860 15934 34862 15986
rect 34862 15934 34914 15986
rect 34914 15934 34916 15986
rect 34860 15932 34916 15934
rect 34636 15202 34692 15204
rect 34636 15150 34638 15202
rect 34638 15150 34690 15202
rect 34690 15150 34692 15202
rect 34636 15148 34692 15150
rect 36204 15932 36260 15988
rect 35644 15820 35700 15876
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 36540 15148 36596 15204
rect 34412 14476 34468 14532
rect 35308 14418 35364 14420
rect 35308 14366 35310 14418
rect 35310 14366 35362 14418
rect 35362 14366 35364 14418
rect 35308 14364 35364 14366
rect 33852 13970 33908 13972
rect 33852 13918 33854 13970
rect 33854 13918 33906 13970
rect 33906 13918 33908 13970
rect 33852 13916 33908 13918
rect 28588 13074 28644 13076
rect 28588 13022 28590 13074
rect 28590 13022 28642 13074
rect 28642 13022 28644 13074
rect 28588 13020 28644 13022
rect 28812 12402 28868 12404
rect 28812 12350 28814 12402
rect 28814 12350 28866 12402
rect 28866 12350 28868 12402
rect 28812 12348 28868 12350
rect 29260 12348 29316 12404
rect 27244 12124 27300 12180
rect 33068 12684 33124 12740
rect 29932 11452 29988 11508
rect 28028 11228 28084 11284
rect 27356 10892 27412 10948
rect 27916 10892 27972 10948
rect 31836 11506 31892 11508
rect 31836 11454 31838 11506
rect 31838 11454 31890 11506
rect 31890 11454 31892 11506
rect 31836 11452 31892 11454
rect 31500 11228 31556 11284
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35868 14530 35924 14532
rect 35868 14478 35870 14530
rect 35870 14478 35922 14530
rect 35922 14478 35924 14530
rect 35868 14476 35924 14478
rect 35644 13132 35700 13188
rect 35532 12684 35588 12740
rect 35868 12738 35924 12740
rect 35868 12686 35870 12738
rect 35870 12686 35922 12738
rect 35922 12686 35924 12738
rect 35868 12684 35924 12686
rect 33964 11900 34020 11956
rect 34972 12348 35028 12404
rect 36092 12738 36148 12740
rect 36092 12686 36094 12738
rect 36094 12686 36146 12738
rect 36146 12686 36148 12738
rect 36092 12684 36148 12686
rect 29820 10892 29876 10948
rect 27020 8428 27076 8484
rect 27580 7586 27636 7588
rect 27580 7534 27582 7586
rect 27582 7534 27634 7586
rect 27634 7534 27636 7586
rect 27580 7532 27636 7534
rect 29372 8876 29428 8932
rect 29036 7980 29092 8036
rect 31500 10108 31556 10164
rect 30268 9996 30324 10052
rect 31164 9436 31220 9492
rect 32508 9772 32564 9828
rect 32732 11228 32788 11284
rect 35980 12178 36036 12180
rect 35980 12126 35982 12178
rect 35982 12126 36034 12178
rect 36034 12126 36036 12178
rect 35980 12124 36036 12126
rect 35196 12066 35252 12068
rect 35196 12014 35198 12066
rect 35198 12014 35250 12066
rect 35250 12014 35252 12066
rect 35196 12012 35252 12014
rect 35420 11900 35476 11956
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 34972 10108 35028 10164
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 34860 9996 34916 10052
rect 36428 12066 36484 12068
rect 36428 12014 36430 12066
rect 36430 12014 36482 12066
rect 36482 12014 36484 12066
rect 36428 12012 36484 12014
rect 36540 11788 36596 11844
rect 35868 9996 35924 10052
rect 32956 9714 33012 9716
rect 32956 9662 32958 9714
rect 32958 9662 33010 9714
rect 33010 9662 33012 9714
rect 32956 9660 33012 9662
rect 30716 8930 30772 8932
rect 30716 8878 30718 8930
rect 30718 8878 30770 8930
rect 30770 8878 30772 8930
rect 30716 8876 30772 8878
rect 30604 8818 30660 8820
rect 30604 8766 30606 8818
rect 30606 8766 30658 8818
rect 30658 8766 30660 8818
rect 30604 8764 30660 8766
rect 29708 7644 29764 7700
rect 26796 6466 26852 6468
rect 26796 6414 26798 6466
rect 26798 6414 26850 6466
rect 26850 6414 26852 6466
rect 26796 6412 26852 6414
rect 27580 6188 27636 6244
rect 27468 6076 27524 6132
rect 28140 5852 28196 5908
rect 26348 4284 26404 4340
rect 29260 5852 29316 5908
rect 30268 7698 30324 7700
rect 30268 7646 30270 7698
rect 30270 7646 30322 7698
rect 30322 7646 30324 7698
rect 30268 7644 30324 7646
rect 30044 7474 30100 7476
rect 30044 7422 30046 7474
rect 30046 7422 30098 7474
rect 30098 7422 30100 7474
rect 30044 7420 30100 7422
rect 29708 5852 29764 5908
rect 28252 5122 28308 5124
rect 28252 5070 28254 5122
rect 28254 5070 28306 5122
rect 28306 5070 28308 5122
rect 28252 5068 28308 5070
rect 29596 5234 29652 5236
rect 29596 5182 29598 5234
rect 29598 5182 29650 5234
rect 29650 5182 29652 5234
rect 29596 5180 29652 5182
rect 30156 5292 30212 5348
rect 31276 8428 31332 8484
rect 33852 9826 33908 9828
rect 33852 9774 33854 9826
rect 33854 9774 33906 9826
rect 33906 9774 33908 9826
rect 33852 9772 33908 9774
rect 35308 9772 35364 9828
rect 33516 9714 33572 9716
rect 33516 9662 33518 9714
rect 33518 9662 33570 9714
rect 33570 9662 33572 9714
rect 33516 9660 33572 9662
rect 33404 8876 33460 8932
rect 35644 9266 35700 9268
rect 35644 9214 35646 9266
rect 35646 9214 35698 9266
rect 35698 9214 35700 9266
rect 35644 9212 35700 9214
rect 35532 8930 35588 8932
rect 35532 8878 35534 8930
rect 35534 8878 35586 8930
rect 35586 8878 35588 8930
rect 35532 8876 35588 8878
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 32284 7644 32340 7700
rect 32172 6802 32228 6804
rect 32172 6750 32174 6802
rect 32174 6750 32226 6802
rect 32226 6750 32228 6802
rect 32172 6748 32228 6750
rect 33180 7698 33236 7700
rect 33180 7646 33182 7698
rect 33182 7646 33234 7698
rect 33234 7646 33236 7698
rect 33180 7644 33236 7646
rect 35980 9714 36036 9716
rect 35980 9662 35982 9714
rect 35982 9662 36034 9714
rect 36034 9662 36036 9714
rect 35980 9660 36036 9662
rect 36204 10332 36260 10388
rect 37548 31276 37604 31332
rect 38108 31500 38164 31556
rect 37772 31106 37828 31108
rect 37772 31054 37774 31106
rect 37774 31054 37826 31106
rect 37826 31054 37828 31106
rect 37772 31052 37828 31054
rect 37884 30994 37940 30996
rect 37884 30942 37886 30994
rect 37886 30942 37938 30994
rect 37938 30942 37940 30994
rect 37884 30940 37940 30942
rect 37996 30044 38052 30100
rect 37548 28812 37604 28868
rect 38220 30268 38276 30324
rect 37660 28700 37716 28756
rect 37884 29650 37940 29652
rect 37884 29598 37886 29650
rect 37886 29598 37938 29650
rect 37938 29598 37940 29650
rect 37884 29596 37940 29598
rect 39452 32450 39508 32452
rect 39452 32398 39454 32450
rect 39454 32398 39506 32450
rect 39506 32398 39508 32450
rect 39452 32396 39508 32398
rect 39116 30994 39172 30996
rect 39116 30942 39118 30994
rect 39118 30942 39170 30994
rect 39170 30942 39172 30994
rect 39116 30940 39172 30942
rect 39228 30770 39284 30772
rect 39228 30718 39230 30770
rect 39230 30718 39282 30770
rect 39282 30718 39284 30770
rect 39228 30716 39284 30718
rect 39004 30268 39060 30324
rect 39452 30044 39508 30100
rect 38444 29596 38500 29652
rect 39004 29650 39060 29652
rect 39004 29598 39006 29650
rect 39006 29598 39058 29650
rect 39058 29598 39060 29650
rect 39004 29596 39060 29598
rect 39788 45612 39844 45668
rect 40236 45836 40292 45892
rect 40572 45836 40628 45892
rect 40236 45666 40292 45668
rect 40236 45614 40238 45666
rect 40238 45614 40290 45666
rect 40290 45614 40292 45666
rect 40236 45612 40292 45614
rect 40012 45052 40068 45108
rect 39676 42642 39732 42644
rect 39676 42590 39678 42642
rect 39678 42590 39730 42642
rect 39730 42590 39732 42642
rect 39676 42588 39732 42590
rect 39900 42588 39956 42644
rect 40348 42754 40404 42756
rect 40348 42702 40350 42754
rect 40350 42702 40402 42754
rect 40402 42702 40404 42754
rect 40348 42700 40404 42702
rect 40236 41020 40292 41076
rect 39788 36988 39844 37044
rect 40012 40402 40068 40404
rect 40012 40350 40014 40402
rect 40014 40350 40066 40402
rect 40066 40350 40068 40402
rect 40012 40348 40068 40350
rect 40236 40348 40292 40404
rect 39900 39676 39956 39732
rect 39676 36652 39732 36708
rect 39788 36258 39844 36260
rect 39788 36206 39790 36258
rect 39790 36206 39842 36258
rect 39842 36206 39844 36258
rect 39788 36204 39844 36206
rect 41132 49196 41188 49252
rect 40908 49026 40964 49028
rect 40908 48974 40910 49026
rect 40910 48974 40962 49026
rect 40962 48974 40964 49026
rect 40908 48972 40964 48974
rect 41356 48914 41412 48916
rect 41356 48862 41358 48914
rect 41358 48862 41410 48914
rect 41410 48862 41412 48914
rect 41356 48860 41412 48862
rect 41020 48130 41076 48132
rect 41020 48078 41022 48130
rect 41022 48078 41074 48130
rect 41074 48078 41076 48130
rect 41020 48076 41076 48078
rect 41580 47458 41636 47460
rect 41580 47406 41582 47458
rect 41582 47406 41634 47458
rect 41634 47406 41636 47458
rect 41580 47404 41636 47406
rect 44156 50428 44212 50484
rect 44940 50482 44996 50484
rect 44940 50430 44942 50482
rect 44942 50430 44994 50482
rect 44994 50430 44996 50482
rect 44940 50428 44996 50430
rect 41804 48130 41860 48132
rect 41804 48078 41806 48130
rect 41806 48078 41858 48130
rect 41858 48078 41860 48130
rect 41804 48076 41860 48078
rect 42476 48076 42532 48132
rect 41916 47346 41972 47348
rect 41916 47294 41918 47346
rect 41918 47294 41970 47346
rect 41970 47294 41972 47346
rect 41916 47292 41972 47294
rect 41804 47234 41860 47236
rect 41804 47182 41806 47234
rect 41806 47182 41858 47234
rect 41858 47182 41860 47234
rect 41804 47180 41860 47182
rect 41132 45836 41188 45892
rect 42700 47346 42756 47348
rect 42700 47294 42702 47346
rect 42702 47294 42754 47346
rect 42754 47294 42756 47346
rect 42700 47292 42756 47294
rect 42924 48076 42980 48132
rect 46396 48802 46452 48804
rect 46396 48750 46398 48802
rect 46398 48750 46450 48802
rect 46450 48750 46452 48802
rect 46396 48748 46452 48750
rect 45500 48076 45556 48132
rect 42476 46620 42532 46676
rect 42252 46396 42308 46452
rect 46172 48130 46228 48132
rect 46172 48078 46174 48130
rect 46174 48078 46226 48130
rect 46226 48078 46228 48130
rect 46172 48076 46228 48078
rect 45724 47180 45780 47236
rect 48300 49698 48356 49700
rect 48300 49646 48302 49698
rect 48302 49646 48354 49698
rect 48354 49646 48356 49698
rect 48300 49644 48356 49646
rect 46956 48802 47012 48804
rect 46956 48750 46958 48802
rect 46958 48750 47010 48802
rect 47010 48750 47012 48802
rect 46956 48748 47012 48750
rect 47180 48914 47236 48916
rect 47180 48862 47182 48914
rect 47182 48862 47234 48914
rect 47234 48862 47236 48914
rect 47180 48860 47236 48862
rect 48748 50370 48804 50372
rect 48748 50318 48750 50370
rect 48750 50318 48802 50370
rect 48802 50318 48804 50370
rect 48748 50316 48804 50318
rect 50652 51378 50708 51380
rect 50652 51326 50654 51378
rect 50654 51326 50706 51378
rect 50706 51326 50708 51378
rect 50652 51324 50708 51326
rect 50428 51212 50484 51268
rect 48748 49026 48804 49028
rect 48748 48974 48750 49026
rect 48750 48974 48802 49026
rect 48802 48974 48804 49026
rect 48748 48972 48804 48974
rect 49196 49698 49252 49700
rect 49196 49646 49198 49698
rect 49198 49646 49250 49698
rect 49250 49646 49252 49698
rect 49196 49644 49252 49646
rect 49980 50316 50036 50372
rect 51212 51378 51268 51380
rect 51212 51326 51214 51378
rect 51214 51326 51266 51378
rect 51266 51326 51268 51378
rect 51212 51324 51268 51326
rect 50556 50202 50612 50204
rect 50556 50150 50558 50202
rect 50558 50150 50610 50202
rect 50610 50150 50612 50202
rect 50556 50148 50612 50150
rect 50660 50202 50716 50204
rect 50660 50150 50662 50202
rect 50662 50150 50714 50202
rect 50714 50150 50716 50202
rect 50660 50148 50716 50150
rect 50764 50202 50820 50204
rect 50764 50150 50766 50202
rect 50766 50150 50818 50202
rect 50818 50150 50820 50202
rect 50764 50148 50820 50150
rect 48412 48860 48468 48916
rect 48972 48860 49028 48916
rect 48188 48748 48244 48804
rect 46844 48242 46900 48244
rect 46844 48190 46846 48242
rect 46846 48190 46898 48242
rect 46898 48190 46900 48242
rect 46844 48188 46900 48190
rect 46732 47292 46788 47348
rect 47180 48076 47236 48132
rect 44156 46508 44212 46564
rect 42924 46396 42980 46452
rect 42028 45890 42084 45892
rect 42028 45838 42030 45890
rect 42030 45838 42082 45890
rect 42082 45838 42084 45890
rect 42028 45836 42084 45838
rect 41468 45724 41524 45780
rect 40908 45106 40964 45108
rect 40908 45054 40910 45106
rect 40910 45054 40962 45106
rect 40962 45054 40964 45106
rect 40908 45052 40964 45054
rect 42364 45778 42420 45780
rect 42364 45726 42366 45778
rect 42366 45726 42418 45778
rect 42418 45726 42420 45778
rect 42364 45724 42420 45726
rect 42252 45276 42308 45332
rect 44380 46396 44436 46452
rect 43260 45890 43316 45892
rect 43260 45838 43262 45890
rect 43262 45838 43314 45890
rect 43314 45838 43316 45890
rect 43260 45836 43316 45838
rect 43148 45778 43204 45780
rect 43148 45726 43150 45778
rect 43150 45726 43202 45778
rect 43202 45726 43204 45778
rect 43148 45724 43204 45726
rect 42924 45666 42980 45668
rect 42924 45614 42926 45666
rect 42926 45614 42978 45666
rect 42978 45614 42980 45666
rect 42924 45612 42980 45614
rect 42700 45500 42756 45556
rect 43148 45500 43204 45556
rect 43820 45778 43876 45780
rect 43820 45726 43822 45778
rect 43822 45726 43874 45778
rect 43874 45726 43876 45778
rect 43820 45724 43876 45726
rect 44044 45500 44100 45556
rect 43372 45276 43428 45332
rect 43260 44994 43316 44996
rect 43260 44942 43262 44994
rect 43262 44942 43314 44994
rect 43314 44942 43316 44994
rect 43260 44940 43316 44942
rect 41356 42812 41412 42868
rect 43148 42866 43204 42868
rect 43148 42814 43150 42866
rect 43150 42814 43202 42866
rect 43202 42814 43204 42866
rect 43148 42812 43204 42814
rect 43820 42700 43876 42756
rect 43932 42812 43988 42868
rect 43484 42642 43540 42644
rect 43484 42590 43486 42642
rect 43486 42590 43538 42642
rect 43538 42590 43540 42642
rect 43484 42588 43540 42590
rect 44268 42754 44324 42756
rect 44268 42702 44270 42754
rect 44270 42702 44322 42754
rect 44322 42702 44324 42754
rect 44268 42700 44324 42702
rect 44492 44994 44548 44996
rect 44492 44942 44494 44994
rect 44494 44942 44546 44994
rect 44546 44942 44548 44994
rect 44492 44940 44548 44942
rect 44828 42812 44884 42868
rect 45388 42812 45444 42868
rect 46060 45276 46116 45332
rect 45948 42812 46004 42868
rect 44268 41804 44324 41860
rect 40348 39564 40404 39620
rect 41132 41020 41188 41076
rect 40348 37154 40404 37156
rect 40348 37102 40350 37154
rect 40350 37102 40402 37154
rect 40402 37102 40404 37154
rect 40348 37100 40404 37102
rect 40012 36204 40068 36260
rect 40796 40402 40852 40404
rect 40796 40350 40798 40402
rect 40798 40350 40850 40402
rect 40850 40350 40852 40402
rect 40796 40348 40852 40350
rect 40908 39340 40964 39396
rect 42028 40626 42084 40628
rect 42028 40574 42030 40626
rect 42030 40574 42082 40626
rect 42082 40574 42084 40626
rect 42028 40572 42084 40574
rect 42364 40236 42420 40292
rect 41468 39788 41524 39844
rect 43036 39788 43092 39844
rect 41356 39618 41412 39620
rect 41356 39566 41358 39618
rect 41358 39566 41410 39618
rect 41410 39566 41412 39618
rect 41356 39564 41412 39566
rect 43036 39004 43092 39060
rect 40908 37996 40964 38052
rect 42812 38722 42868 38724
rect 42812 38670 42814 38722
rect 42814 38670 42866 38722
rect 42866 38670 42868 38722
rect 42812 38668 42868 38670
rect 40460 36092 40516 36148
rect 40908 35532 40964 35588
rect 39900 34130 39956 34132
rect 39900 34078 39902 34130
rect 39902 34078 39954 34130
rect 39954 34078 39956 34130
rect 39900 34076 39956 34078
rect 39676 31778 39732 31780
rect 39676 31726 39678 31778
rect 39678 31726 39730 31778
rect 39730 31726 39732 31778
rect 39676 31724 39732 31726
rect 39676 29484 39732 29540
rect 39004 29426 39060 29428
rect 39004 29374 39006 29426
rect 39006 29374 39058 29426
rect 39058 29374 39060 29426
rect 39004 29372 39060 29374
rect 38220 29148 38276 29204
rect 39564 29260 39620 29316
rect 39340 29202 39396 29204
rect 39340 29150 39342 29202
rect 39342 29150 39394 29202
rect 39394 29150 39396 29202
rect 39340 29148 39396 29150
rect 39004 28812 39060 28868
rect 37436 28028 37492 28084
rect 37660 27858 37716 27860
rect 37660 27806 37662 27858
rect 37662 27806 37714 27858
rect 37714 27806 37716 27858
rect 37660 27804 37716 27806
rect 37212 27746 37268 27748
rect 37212 27694 37214 27746
rect 37214 27694 37266 27746
rect 37266 27694 37268 27746
rect 37212 27692 37268 27694
rect 37772 27020 37828 27076
rect 37884 27916 37940 27972
rect 37324 26124 37380 26180
rect 37100 25452 37156 25508
rect 36988 24108 37044 24164
rect 37100 24722 37156 24724
rect 37100 24670 37102 24722
rect 37102 24670 37154 24722
rect 37154 24670 37156 24722
rect 37100 24668 37156 24670
rect 36988 22370 37044 22372
rect 36988 22318 36990 22370
rect 36990 22318 37042 22370
rect 37042 22318 37044 22370
rect 36988 22316 37044 22318
rect 37548 25282 37604 25284
rect 37548 25230 37550 25282
rect 37550 25230 37602 25282
rect 37602 25230 37604 25282
rect 37548 25228 37604 25230
rect 37660 25004 37716 25060
rect 37772 24722 37828 24724
rect 37772 24670 37774 24722
rect 37774 24670 37826 24722
rect 37826 24670 37828 24722
rect 37772 24668 37828 24670
rect 37660 23938 37716 23940
rect 37660 23886 37662 23938
rect 37662 23886 37714 23938
rect 37714 23886 37716 23938
rect 37660 23884 37716 23886
rect 37324 23660 37380 23716
rect 37212 23042 37268 23044
rect 37212 22990 37214 23042
rect 37214 22990 37266 23042
rect 37266 22990 37268 23042
rect 37212 22988 37268 22990
rect 37324 22258 37380 22260
rect 37324 22206 37326 22258
rect 37326 22206 37378 22258
rect 37378 22206 37380 22258
rect 37324 22204 37380 22206
rect 37212 21756 37268 21812
rect 37100 21420 37156 21476
rect 36764 16716 36820 16772
rect 37100 15372 37156 15428
rect 36988 15314 37044 15316
rect 36988 15262 36990 15314
rect 36990 15262 37042 15314
rect 37042 15262 37044 15314
rect 36988 15260 37044 15262
rect 37100 12178 37156 12180
rect 37100 12126 37102 12178
rect 37102 12126 37154 12178
rect 37154 12126 37156 12178
rect 37100 12124 37156 12126
rect 37548 22988 37604 23044
rect 37548 21868 37604 21924
rect 39900 32674 39956 32676
rect 39900 32622 39902 32674
rect 39902 32622 39954 32674
rect 39954 32622 39956 32674
rect 39900 32620 39956 32622
rect 40236 35308 40292 35364
rect 39900 31778 39956 31780
rect 39900 31726 39902 31778
rect 39902 31726 39954 31778
rect 39954 31726 39956 31778
rect 39900 31724 39956 31726
rect 40796 34860 40852 34916
rect 42364 37324 42420 37380
rect 42028 36988 42084 37044
rect 41020 33404 41076 33460
rect 40460 32674 40516 32676
rect 40460 32622 40462 32674
rect 40462 32622 40514 32674
rect 40514 32622 40516 32674
rect 40460 32620 40516 32622
rect 40236 31948 40292 32004
rect 40908 31948 40964 32004
rect 40348 31724 40404 31780
rect 40348 29538 40404 29540
rect 40348 29486 40350 29538
rect 40350 29486 40402 29538
rect 40402 29486 40404 29538
rect 40348 29484 40404 29486
rect 41020 31724 41076 31780
rect 41468 34860 41524 34916
rect 41916 34690 41972 34692
rect 41916 34638 41918 34690
rect 41918 34638 41970 34690
rect 41970 34638 41972 34690
rect 41916 34636 41972 34638
rect 44940 41804 44996 41860
rect 44268 41020 44324 41076
rect 43708 40514 43764 40516
rect 43708 40462 43710 40514
rect 43710 40462 43762 40514
rect 43762 40462 43764 40514
rect 43708 40460 43764 40462
rect 44492 40460 44548 40516
rect 43932 40236 43988 40292
rect 44268 39452 44324 39508
rect 43932 38668 43988 38724
rect 42812 34972 42868 35028
rect 42140 34076 42196 34132
rect 41468 33404 41524 33460
rect 41804 33404 41860 33460
rect 40684 29372 40740 29428
rect 40236 28252 40292 28308
rect 39788 27580 39844 27636
rect 39788 27186 39844 27188
rect 39788 27134 39790 27186
rect 39790 27134 39842 27186
rect 39842 27134 39844 27186
rect 39788 27132 39844 27134
rect 37996 26796 38052 26852
rect 37996 25788 38052 25844
rect 39900 26908 39956 26964
rect 39452 26684 39508 26740
rect 38780 26290 38836 26292
rect 38780 26238 38782 26290
rect 38782 26238 38834 26290
rect 38834 26238 38836 26290
rect 38780 26236 38836 26238
rect 38892 26066 38948 26068
rect 38892 26014 38894 26066
rect 38894 26014 38946 26066
rect 38946 26014 38948 26066
rect 38892 26012 38948 26014
rect 39676 26012 39732 26068
rect 38668 25676 38724 25732
rect 39340 25788 39396 25844
rect 38108 25452 38164 25508
rect 37996 23826 38052 23828
rect 37996 23774 37998 23826
rect 37998 23774 38050 23826
rect 38050 23774 38052 23826
rect 37996 23772 38052 23774
rect 38556 25282 38612 25284
rect 38556 25230 38558 25282
rect 38558 25230 38610 25282
rect 38610 25230 38612 25282
rect 38556 25228 38612 25230
rect 38556 24722 38612 24724
rect 38556 24670 38558 24722
rect 38558 24670 38610 24722
rect 38610 24670 38612 24722
rect 38556 24668 38612 24670
rect 38780 23826 38836 23828
rect 38780 23774 38782 23826
rect 38782 23774 38834 23826
rect 38834 23774 38836 23826
rect 38780 23772 38836 23774
rect 38444 22988 38500 23044
rect 38556 21810 38612 21812
rect 38556 21758 38558 21810
rect 38558 21758 38610 21810
rect 38610 21758 38612 21810
rect 38556 21756 38612 21758
rect 37996 21644 38052 21700
rect 37660 21420 37716 21476
rect 38108 21474 38164 21476
rect 38108 21422 38110 21474
rect 38110 21422 38162 21474
rect 38162 21422 38164 21474
rect 38108 21420 38164 21422
rect 37548 20860 37604 20916
rect 39340 25394 39396 25396
rect 39340 25342 39342 25394
rect 39342 25342 39394 25394
rect 39394 25342 39396 25394
rect 39340 25340 39396 25342
rect 39452 24892 39508 24948
rect 39788 24892 39844 24948
rect 39900 25340 39956 25396
rect 40124 26684 40180 26740
rect 39676 24556 39732 24612
rect 39564 23884 39620 23940
rect 39452 23436 39508 23492
rect 39228 22316 39284 22372
rect 39228 21644 39284 21700
rect 39564 20524 39620 20580
rect 39004 19628 39060 19684
rect 40012 24444 40068 24500
rect 39788 19794 39844 19796
rect 39788 19742 39790 19794
rect 39790 19742 39842 19794
rect 39842 19742 39844 19794
rect 39788 19740 39844 19742
rect 39788 19516 39844 19572
rect 38444 19458 38500 19460
rect 38444 19406 38446 19458
rect 38446 19406 38498 19458
rect 38498 19406 38500 19458
rect 38444 19404 38500 19406
rect 38332 18508 38388 18564
rect 38892 18450 38948 18452
rect 38892 18398 38894 18450
rect 38894 18398 38946 18450
rect 38946 18398 38948 18450
rect 38892 18396 38948 18398
rect 38556 17724 38612 17780
rect 37884 17388 37940 17444
rect 37436 10892 37492 10948
rect 38108 17666 38164 17668
rect 38108 17614 38110 17666
rect 38110 17614 38162 17666
rect 38162 17614 38164 17666
rect 38108 17612 38164 17614
rect 38556 17554 38612 17556
rect 38556 17502 38558 17554
rect 38558 17502 38610 17554
rect 38610 17502 38612 17554
rect 38556 17500 38612 17502
rect 37772 15874 37828 15876
rect 37772 15822 37774 15874
rect 37774 15822 37826 15874
rect 37826 15822 37828 15874
rect 37772 15820 37828 15822
rect 38108 15932 38164 15988
rect 38220 16380 38276 16436
rect 38668 16268 38724 16324
rect 38556 16156 38612 16212
rect 37996 15820 38052 15876
rect 40012 23154 40068 23156
rect 40012 23102 40014 23154
rect 40014 23102 40066 23154
rect 40066 23102 40068 23154
rect 40012 23100 40068 23102
rect 40012 22316 40068 22372
rect 40236 25116 40292 25172
rect 40348 21644 40404 21700
rect 40460 22092 40516 22148
rect 40124 20188 40180 20244
rect 40236 21586 40292 21588
rect 40236 21534 40238 21586
rect 40238 21534 40290 21586
rect 40290 21534 40292 21586
rect 40236 21532 40292 21534
rect 40348 18396 40404 18452
rect 39452 16380 39508 16436
rect 39564 17724 39620 17780
rect 38668 15596 38724 15652
rect 38332 15148 38388 15204
rect 38444 15372 38500 15428
rect 39564 15484 39620 15540
rect 38780 14924 38836 14980
rect 38892 14588 38948 14644
rect 38108 14364 38164 14420
rect 38108 13132 38164 13188
rect 38332 12962 38388 12964
rect 38332 12910 38334 12962
rect 38334 12910 38386 12962
rect 38386 12910 38388 12962
rect 38332 12908 38388 12910
rect 39228 13244 39284 13300
rect 37772 12684 37828 12740
rect 38220 11788 38276 11844
rect 38556 12738 38612 12740
rect 38556 12686 38558 12738
rect 38558 12686 38610 12738
rect 38610 12686 38612 12738
rect 38556 12684 38612 12686
rect 39788 15426 39844 15428
rect 39788 15374 39790 15426
rect 39790 15374 39842 15426
rect 39842 15374 39844 15426
rect 39788 15372 39844 15374
rect 39676 14252 39732 14308
rect 37660 9996 37716 10052
rect 38220 9826 38276 9828
rect 38220 9774 38222 9826
rect 38222 9774 38274 9826
rect 38274 9774 38276 9826
rect 38220 9772 38276 9774
rect 38668 9826 38724 9828
rect 38668 9774 38670 9826
rect 38670 9774 38722 9826
rect 38722 9774 38724 9826
rect 38668 9772 38724 9774
rect 39900 14924 39956 14980
rect 40236 14924 40292 14980
rect 40012 14140 40068 14196
rect 40012 12908 40068 12964
rect 39676 9772 39732 9828
rect 37100 9548 37156 9604
rect 35756 7420 35812 7476
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 33292 6860 33348 6916
rect 31724 6076 31780 6132
rect 32508 6524 32564 6580
rect 31500 5346 31556 5348
rect 31500 5294 31502 5346
rect 31502 5294 31554 5346
rect 31554 5294 31556 5346
rect 31500 5292 31556 5294
rect 30380 5180 30436 5236
rect 33068 6130 33124 6132
rect 33068 6078 33070 6130
rect 33070 6078 33122 6130
rect 33122 6078 33124 6130
rect 33068 6076 33124 6078
rect 33628 6578 33684 6580
rect 33628 6526 33630 6578
rect 33630 6526 33682 6578
rect 33682 6526 33684 6578
rect 33628 6524 33684 6526
rect 36204 6802 36260 6804
rect 36204 6750 36206 6802
rect 36206 6750 36258 6802
rect 36258 6750 36260 6802
rect 36204 6748 36260 6750
rect 37660 9548 37716 9604
rect 37996 9212 38052 9268
rect 37324 8204 37380 8260
rect 37548 7532 37604 7588
rect 37436 6524 37492 6580
rect 33740 5906 33796 5908
rect 33740 5854 33742 5906
rect 33742 5854 33794 5906
rect 33794 5854 33796 5906
rect 33740 5852 33796 5854
rect 37996 8034 38052 8036
rect 37996 7982 37998 8034
rect 37998 7982 38050 8034
rect 38050 7982 38052 8034
rect 37996 7980 38052 7982
rect 38332 7756 38388 7812
rect 38780 7308 38836 7364
rect 38220 6690 38276 6692
rect 38220 6638 38222 6690
rect 38222 6638 38274 6690
rect 38274 6638 38276 6690
rect 38220 6636 38276 6638
rect 38780 6636 38836 6692
rect 38332 6524 38388 6580
rect 39228 9548 39284 9604
rect 39788 12684 39844 12740
rect 39564 7980 39620 8036
rect 39228 6578 39284 6580
rect 39228 6526 39230 6578
rect 39230 6526 39282 6578
rect 39282 6526 39284 6578
rect 39228 6524 39284 6526
rect 35980 5906 36036 5908
rect 35980 5854 35982 5906
rect 35982 5854 36034 5906
rect 36034 5854 36036 5906
rect 35980 5852 36036 5854
rect 36204 5852 36260 5908
rect 32956 5180 33012 5236
rect 28364 5010 28420 5012
rect 28364 4958 28366 5010
rect 28366 4958 28418 5010
rect 28418 4958 28420 5010
rect 28364 4956 28420 4958
rect 31612 4956 31668 5012
rect 32172 4956 32228 5012
rect 28812 4226 28868 4228
rect 28812 4174 28814 4226
rect 28814 4174 28866 4226
rect 28866 4174 28868 4226
rect 28812 4172 28868 4174
rect 29260 4338 29316 4340
rect 29260 4286 29262 4338
rect 29262 4286 29314 4338
rect 29314 4286 29316 4338
rect 29260 4284 29316 4286
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 36428 5234 36484 5236
rect 36428 5182 36430 5234
rect 36430 5182 36482 5234
rect 36482 5182 36484 5234
rect 36428 5180 36484 5182
rect 36876 5180 36932 5236
rect 37212 5906 37268 5908
rect 37212 5854 37214 5906
rect 37214 5854 37266 5906
rect 37266 5854 37268 5906
rect 37212 5852 37268 5854
rect 41804 32956 41860 33012
rect 40908 30268 40964 30324
rect 41132 29986 41188 29988
rect 41132 29934 41134 29986
rect 41134 29934 41186 29986
rect 41186 29934 41188 29986
rect 41132 29932 41188 29934
rect 42028 29986 42084 29988
rect 42028 29934 42030 29986
rect 42030 29934 42082 29986
rect 42082 29934 42084 29986
rect 42028 29932 42084 29934
rect 42700 34076 42756 34132
rect 44044 37378 44100 37380
rect 44044 37326 44046 37378
rect 44046 37326 44098 37378
rect 44098 37326 44100 37378
rect 44044 37324 44100 37326
rect 43484 35756 43540 35812
rect 44044 36316 44100 36372
rect 43932 34972 43988 35028
rect 43148 34636 43204 34692
rect 42476 33516 42532 33572
rect 43372 33516 43428 33572
rect 43372 32956 43428 33012
rect 44492 35810 44548 35812
rect 44492 35758 44494 35810
rect 44494 35758 44546 35810
rect 44546 35758 44548 35810
rect 44492 35756 44548 35758
rect 44828 34972 44884 35028
rect 45276 41858 45332 41860
rect 45276 41806 45278 41858
rect 45278 41806 45330 41858
rect 45330 41806 45332 41858
rect 45276 41804 45332 41806
rect 45836 41074 45892 41076
rect 45836 41022 45838 41074
rect 45838 41022 45890 41074
rect 45890 41022 45892 41074
rect 45836 41020 45892 41022
rect 45724 40962 45780 40964
rect 45724 40910 45726 40962
rect 45726 40910 45778 40962
rect 45778 40910 45780 40962
rect 45724 40908 45780 40910
rect 48188 47964 48244 48020
rect 46508 46562 46564 46564
rect 46508 46510 46510 46562
rect 46510 46510 46562 46562
rect 46562 46510 46564 46562
rect 46508 46508 46564 46510
rect 46620 45276 46676 45332
rect 48188 46674 48244 46676
rect 48188 46622 48190 46674
rect 48190 46622 48242 46674
rect 48242 46622 48244 46674
rect 48188 46620 48244 46622
rect 49308 48188 49364 48244
rect 48748 47346 48804 47348
rect 48748 47294 48750 47346
rect 48750 47294 48802 47346
rect 48802 47294 48804 47346
rect 48748 47292 48804 47294
rect 48972 48018 49028 48020
rect 48972 47966 48974 48018
rect 48974 47966 49026 48018
rect 49026 47966 49028 48018
rect 48972 47964 49028 47966
rect 48860 46844 48916 46900
rect 48748 46674 48804 46676
rect 48748 46622 48750 46674
rect 48750 46622 48802 46674
rect 48802 46622 48804 46674
rect 48748 46620 48804 46622
rect 49308 46562 49364 46564
rect 49308 46510 49310 46562
rect 49310 46510 49362 46562
rect 49362 46510 49364 46562
rect 49308 46508 49364 46510
rect 49308 45836 49364 45892
rect 48748 45164 48804 45220
rect 49980 48972 50036 49028
rect 49980 48188 50036 48244
rect 49868 47292 49924 47348
rect 50204 49196 50260 49252
rect 51436 51212 51492 51268
rect 50428 49196 50484 49252
rect 50556 48634 50612 48636
rect 50556 48582 50558 48634
rect 50558 48582 50610 48634
rect 50610 48582 50612 48634
rect 50556 48580 50612 48582
rect 50660 48634 50716 48636
rect 50660 48582 50662 48634
rect 50662 48582 50714 48634
rect 50714 48582 50716 48634
rect 50660 48580 50716 48582
rect 50764 48634 50820 48636
rect 50764 48582 50766 48634
rect 50766 48582 50818 48634
rect 50818 48582 50820 48634
rect 50764 48580 50820 48582
rect 50556 47066 50612 47068
rect 50556 47014 50558 47066
rect 50558 47014 50610 47066
rect 50610 47014 50612 47066
rect 50556 47012 50612 47014
rect 50660 47066 50716 47068
rect 50660 47014 50662 47066
rect 50662 47014 50714 47066
rect 50714 47014 50716 47066
rect 50660 47012 50716 47014
rect 50764 47066 50820 47068
rect 50764 47014 50766 47066
rect 50766 47014 50818 47066
rect 50818 47014 50820 47066
rect 50764 47012 50820 47014
rect 53228 49084 53284 49140
rect 51884 48860 51940 48916
rect 50988 46620 51044 46676
rect 48300 45052 48356 45108
rect 47516 43484 47572 43540
rect 46956 42700 47012 42756
rect 46956 41916 47012 41972
rect 47180 43372 47236 43428
rect 45276 39340 45332 39396
rect 45276 36428 45332 36484
rect 43708 34130 43764 34132
rect 43708 34078 43710 34130
rect 43710 34078 43762 34130
rect 43762 34078 43764 34130
rect 43708 34076 43764 34078
rect 43596 32786 43652 32788
rect 43596 32734 43598 32786
rect 43598 32734 43650 32786
rect 43650 32734 43652 32786
rect 43596 32732 43652 32734
rect 42588 32284 42644 32340
rect 43148 32284 43204 32340
rect 42924 32172 42980 32228
rect 42252 31612 42308 31668
rect 42028 29708 42084 29764
rect 41244 29538 41300 29540
rect 41244 29486 41246 29538
rect 41246 29486 41298 29538
rect 41298 29486 41300 29538
rect 41244 29484 41300 29486
rect 41132 28700 41188 28756
rect 41356 28082 41412 28084
rect 41356 28030 41358 28082
rect 41358 28030 41410 28082
rect 41410 28030 41412 28082
rect 41356 28028 41412 28030
rect 41356 27244 41412 27300
rect 41468 27074 41524 27076
rect 41468 27022 41470 27074
rect 41470 27022 41522 27074
rect 41522 27022 41524 27074
rect 41468 27020 41524 27022
rect 42140 29538 42196 29540
rect 42140 29486 42142 29538
rect 42142 29486 42194 29538
rect 42194 29486 42196 29538
rect 42140 29484 42196 29486
rect 41916 28700 41972 28756
rect 42812 31778 42868 31780
rect 42812 31726 42814 31778
rect 42814 31726 42866 31778
rect 42866 31726 42868 31778
rect 42812 31724 42868 31726
rect 43372 31724 43428 31780
rect 43932 32956 43988 33012
rect 43596 32060 43652 32116
rect 42700 31666 42756 31668
rect 42700 31614 42702 31666
rect 42702 31614 42754 31666
rect 42754 31614 42756 31666
rect 42700 31612 42756 31614
rect 42812 31388 42868 31444
rect 43372 31388 43428 31444
rect 43036 30994 43092 30996
rect 43036 30942 43038 30994
rect 43038 30942 43090 30994
rect 43090 30942 43092 30994
rect 43036 30940 43092 30942
rect 42588 30210 42644 30212
rect 42588 30158 42590 30210
rect 42590 30158 42642 30210
rect 42642 30158 42644 30210
rect 42588 30156 42644 30158
rect 42588 29708 42644 29764
rect 42924 28866 42980 28868
rect 42924 28814 42926 28866
rect 42926 28814 42978 28866
rect 42978 28814 42980 28866
rect 42924 28812 42980 28814
rect 43708 31724 43764 31780
rect 43820 31388 43876 31444
rect 43820 31218 43876 31220
rect 43820 31166 43822 31218
rect 43822 31166 43874 31218
rect 43874 31166 43876 31218
rect 43820 31164 43876 31166
rect 43708 31106 43764 31108
rect 43708 31054 43710 31106
rect 43710 31054 43762 31106
rect 43762 31054 43764 31106
rect 43708 31052 43764 31054
rect 43484 28754 43540 28756
rect 43484 28702 43486 28754
rect 43486 28702 43538 28754
rect 43538 28702 43540 28754
rect 43484 28700 43540 28702
rect 42924 28642 42980 28644
rect 42924 28590 42926 28642
rect 42926 28590 42978 28642
rect 42978 28590 42980 28642
rect 42924 28588 42980 28590
rect 43260 28364 43316 28420
rect 43372 28476 43428 28532
rect 41804 28028 41860 28084
rect 45612 39564 45668 39620
rect 46060 39506 46116 39508
rect 46060 39454 46062 39506
rect 46062 39454 46114 39506
rect 46114 39454 46116 39506
rect 46060 39452 46116 39454
rect 46284 39564 46340 39620
rect 45724 38834 45780 38836
rect 45724 38782 45726 38834
rect 45726 38782 45778 38834
rect 45778 38782 45780 38834
rect 45724 38780 45780 38782
rect 46844 39564 46900 39620
rect 46396 39058 46452 39060
rect 46396 39006 46398 39058
rect 46398 39006 46450 39058
rect 46450 39006 46452 39058
rect 46396 39004 46452 39006
rect 46284 38780 46340 38836
rect 46956 39116 47012 39172
rect 48300 43426 48356 43428
rect 48300 43374 48302 43426
rect 48302 43374 48354 43426
rect 48354 43374 48356 43426
rect 48300 43372 48356 43374
rect 48748 42924 48804 42980
rect 48972 45106 49028 45108
rect 48972 45054 48974 45106
rect 48974 45054 49026 45106
rect 49026 45054 49028 45106
rect 48972 45052 49028 45054
rect 50204 45836 50260 45892
rect 49196 45666 49252 45668
rect 49196 45614 49198 45666
rect 49198 45614 49250 45666
rect 49250 45614 49252 45666
rect 49196 45612 49252 45614
rect 49084 44604 49140 44660
rect 48972 43372 49028 43428
rect 49868 45612 49924 45668
rect 50092 45218 50148 45220
rect 50092 45166 50094 45218
rect 50094 45166 50146 45218
rect 50146 45166 50148 45218
rect 50092 45164 50148 45166
rect 49756 44604 49812 44660
rect 49644 44156 49700 44212
rect 49196 43372 49252 43428
rect 48076 41970 48132 41972
rect 48076 41918 48078 41970
rect 48078 41918 48130 41970
rect 48130 41918 48132 41970
rect 48076 41916 48132 41918
rect 47404 40908 47460 40964
rect 47292 39004 47348 39060
rect 46172 36482 46228 36484
rect 46172 36430 46174 36482
rect 46174 36430 46226 36482
rect 46226 36430 46228 36482
rect 46172 36428 46228 36430
rect 46956 37100 47012 37156
rect 46060 36316 46116 36372
rect 46284 35698 46340 35700
rect 46284 35646 46286 35698
rect 46286 35646 46338 35698
rect 46338 35646 46340 35698
rect 46284 35644 46340 35646
rect 45948 35308 46004 35364
rect 45500 34300 45556 34356
rect 45948 33628 46004 33684
rect 45612 33346 45668 33348
rect 45612 33294 45614 33346
rect 45614 33294 45666 33346
rect 45666 33294 45668 33346
rect 45612 33292 45668 33294
rect 45164 32060 45220 32116
rect 44156 31778 44212 31780
rect 44156 31726 44158 31778
rect 44158 31726 44210 31778
rect 44210 31726 44212 31778
rect 44156 31724 44212 31726
rect 44380 31500 44436 31556
rect 44044 31106 44100 31108
rect 44044 31054 44046 31106
rect 44046 31054 44098 31106
rect 44098 31054 44100 31106
rect 44044 31052 44100 31054
rect 44828 31106 44884 31108
rect 44828 31054 44830 31106
rect 44830 31054 44882 31106
rect 44882 31054 44884 31106
rect 44828 31052 44884 31054
rect 44604 28588 44660 28644
rect 43708 27746 43764 27748
rect 43708 27694 43710 27746
rect 43710 27694 43762 27746
rect 43762 27694 43764 27746
rect 43708 27692 43764 27694
rect 42028 26908 42084 26964
rect 40796 25340 40852 25396
rect 40908 21868 40964 21924
rect 41356 26124 41412 26180
rect 41244 24556 41300 24612
rect 41356 22764 41412 22820
rect 41244 22370 41300 22372
rect 41244 22318 41246 22370
rect 41246 22318 41298 22370
rect 41298 22318 41300 22370
rect 41244 22316 41300 22318
rect 43036 27020 43092 27076
rect 42364 26514 42420 26516
rect 42364 26462 42366 26514
rect 42366 26462 42418 26514
rect 42418 26462 42420 26514
rect 42364 26460 42420 26462
rect 42140 26124 42196 26180
rect 42924 26178 42980 26180
rect 42924 26126 42926 26178
rect 42926 26126 42978 26178
rect 42978 26126 42980 26178
rect 42924 26124 42980 26126
rect 42252 25282 42308 25284
rect 42252 25230 42254 25282
rect 42254 25230 42306 25282
rect 42306 25230 42308 25282
rect 42252 25228 42308 25230
rect 42252 24722 42308 24724
rect 42252 24670 42254 24722
rect 42254 24670 42306 24722
rect 42306 24670 42308 24722
rect 42252 24668 42308 24670
rect 42140 24444 42196 24500
rect 42140 23042 42196 23044
rect 42140 22990 42142 23042
rect 42142 22990 42194 23042
rect 42194 22990 42196 23042
rect 42140 22988 42196 22990
rect 41468 22204 41524 22260
rect 41692 22092 41748 22148
rect 41356 21868 41412 21924
rect 41580 21644 41636 21700
rect 41132 21586 41188 21588
rect 41132 21534 41134 21586
rect 41134 21534 41186 21586
rect 41186 21534 41188 21586
rect 41132 21532 41188 21534
rect 41244 21362 41300 21364
rect 41244 21310 41246 21362
rect 41246 21310 41298 21362
rect 41298 21310 41300 21362
rect 41244 21308 41300 21310
rect 41020 21084 41076 21140
rect 40908 19906 40964 19908
rect 40908 19854 40910 19906
rect 40910 19854 40962 19906
rect 40962 19854 40964 19906
rect 40908 19852 40964 19854
rect 42588 23436 42644 23492
rect 42700 23042 42756 23044
rect 42700 22990 42702 23042
rect 42702 22990 42754 23042
rect 42754 22990 42756 23042
rect 42700 22988 42756 22990
rect 43708 26908 43764 26964
rect 43148 25004 43204 25060
rect 44156 27074 44212 27076
rect 44156 27022 44158 27074
rect 44158 27022 44210 27074
rect 44210 27022 44212 27074
rect 44156 27020 44212 27022
rect 42924 22988 42980 23044
rect 42588 22930 42644 22932
rect 42588 22878 42590 22930
rect 42590 22878 42642 22930
rect 42642 22878 42644 22930
rect 42588 22876 42644 22878
rect 42364 22092 42420 22148
rect 42700 22370 42756 22372
rect 42700 22318 42702 22370
rect 42702 22318 42754 22370
rect 42754 22318 42756 22370
rect 42700 22316 42756 22318
rect 42700 22092 42756 22148
rect 42812 21756 42868 21812
rect 43036 21644 43092 21700
rect 43148 24610 43204 24612
rect 43148 24558 43150 24610
rect 43150 24558 43202 24610
rect 43202 24558 43204 24610
rect 43148 24556 43204 24558
rect 42812 21308 42868 21364
rect 42140 18844 42196 18900
rect 44044 25004 44100 25060
rect 43484 24722 43540 24724
rect 43484 24670 43486 24722
rect 43486 24670 43538 24722
rect 43538 24670 43540 24722
rect 43484 24668 43540 24670
rect 43596 23826 43652 23828
rect 43596 23774 43598 23826
rect 43598 23774 43650 23826
rect 43650 23774 43652 23826
rect 43596 23772 43652 23774
rect 43260 23324 43316 23380
rect 43484 23100 43540 23156
rect 43260 22764 43316 22820
rect 43484 22316 43540 22372
rect 43596 23436 43652 23492
rect 43820 22146 43876 22148
rect 43820 22094 43822 22146
rect 43822 22094 43874 22146
rect 43874 22094 43876 22146
rect 43820 22092 43876 22094
rect 44044 23826 44100 23828
rect 44044 23774 44046 23826
rect 44046 23774 44098 23826
rect 44098 23774 44100 23826
rect 44044 23772 44100 23774
rect 44156 23154 44212 23156
rect 44156 23102 44158 23154
rect 44158 23102 44210 23154
rect 44210 23102 44212 23154
rect 44156 23100 44212 23102
rect 44268 22146 44324 22148
rect 44268 22094 44270 22146
rect 44270 22094 44322 22146
rect 44322 22094 44324 22146
rect 44268 22092 44324 22094
rect 43596 21810 43652 21812
rect 43596 21758 43598 21810
rect 43598 21758 43650 21810
rect 43650 21758 43652 21810
rect 43596 21756 43652 21758
rect 43484 21644 43540 21700
rect 43932 21586 43988 21588
rect 43932 21534 43934 21586
rect 43934 21534 43986 21586
rect 43986 21534 43988 21586
rect 43932 21532 43988 21534
rect 45164 31500 45220 31556
rect 45164 30940 45220 30996
rect 44940 29596 44996 29652
rect 45052 28588 45108 28644
rect 45276 27692 45332 27748
rect 45612 32396 45668 32452
rect 48188 36988 48244 37044
rect 47292 30156 47348 30212
rect 47404 34636 47460 34692
rect 47068 30044 47124 30100
rect 46508 28754 46564 28756
rect 46508 28702 46510 28754
rect 46510 28702 46562 28754
rect 46562 28702 46564 28754
rect 46508 28700 46564 28702
rect 45500 27746 45556 27748
rect 45500 27694 45502 27746
rect 45502 27694 45554 27746
rect 45554 27694 45556 27746
rect 45500 27692 45556 27694
rect 45500 27132 45556 27188
rect 46060 25506 46116 25508
rect 46060 25454 46062 25506
rect 46062 25454 46114 25506
rect 46114 25454 46116 25506
rect 46060 25452 46116 25454
rect 44604 23548 44660 23604
rect 44828 23772 44884 23828
rect 44492 23042 44548 23044
rect 44492 22990 44494 23042
rect 44494 22990 44546 23042
rect 44546 22990 44548 23042
rect 44492 22988 44548 22990
rect 44492 22092 44548 22148
rect 45388 23436 45444 23492
rect 45724 23548 45780 23604
rect 46172 25340 46228 25396
rect 46396 25116 46452 25172
rect 46172 23938 46228 23940
rect 46172 23886 46174 23938
rect 46174 23886 46226 23938
rect 46226 23886 46228 23938
rect 46172 23884 46228 23886
rect 45612 23324 45668 23380
rect 45052 22146 45108 22148
rect 45052 22094 45054 22146
rect 45054 22094 45106 22146
rect 45106 22094 45108 22146
rect 45052 22092 45108 22094
rect 45388 22258 45444 22260
rect 45388 22206 45390 22258
rect 45390 22206 45442 22258
rect 45442 22206 45444 22258
rect 45388 22204 45444 22206
rect 46396 23324 46452 23380
rect 46284 22876 46340 22932
rect 46284 22204 46340 22260
rect 45388 21868 45444 21924
rect 45276 21532 45332 21588
rect 44940 20690 44996 20692
rect 44940 20638 44942 20690
rect 44942 20638 44994 20690
rect 44994 20638 44996 20690
rect 44940 20636 44996 20638
rect 43260 20188 43316 20244
rect 43372 18844 43428 18900
rect 42028 18508 42084 18564
rect 42588 18508 42644 18564
rect 41020 18396 41076 18452
rect 41804 18450 41860 18452
rect 41804 18398 41806 18450
rect 41806 18398 41858 18450
rect 41858 18398 41860 18450
rect 41804 18396 41860 18398
rect 41916 18284 41972 18340
rect 40460 17666 40516 17668
rect 40460 17614 40462 17666
rect 40462 17614 40514 17666
rect 40514 17614 40516 17666
rect 40460 17612 40516 17614
rect 42252 18450 42308 18452
rect 42252 18398 42254 18450
rect 42254 18398 42306 18450
rect 42306 18398 42308 18450
rect 42252 18396 42308 18398
rect 42028 16940 42084 16996
rect 41020 16156 41076 16212
rect 40796 16098 40852 16100
rect 40796 16046 40798 16098
rect 40798 16046 40850 16098
rect 40850 16046 40852 16098
rect 40796 16044 40852 16046
rect 40684 15986 40740 15988
rect 40684 15934 40686 15986
rect 40686 15934 40738 15986
rect 40738 15934 40740 15986
rect 40684 15932 40740 15934
rect 40348 12348 40404 12404
rect 40460 13244 40516 13300
rect 40684 14588 40740 14644
rect 41468 15820 41524 15876
rect 41244 15314 41300 15316
rect 41244 15262 41246 15314
rect 41246 15262 41298 15314
rect 41298 15262 41300 15314
rect 41244 15260 41300 15262
rect 42924 18338 42980 18340
rect 42924 18286 42926 18338
rect 42926 18286 42978 18338
rect 42978 18286 42980 18338
rect 42924 18284 42980 18286
rect 43260 18284 43316 18340
rect 42700 16994 42756 16996
rect 42700 16942 42702 16994
rect 42702 16942 42754 16994
rect 42754 16942 42756 16994
rect 42700 16940 42756 16942
rect 42364 15426 42420 15428
rect 42364 15374 42366 15426
rect 42366 15374 42418 15426
rect 42418 15374 42420 15426
rect 42364 15372 42420 15374
rect 42476 15314 42532 15316
rect 42476 15262 42478 15314
rect 42478 15262 42530 15314
rect 42530 15262 42532 15314
rect 42476 15260 42532 15262
rect 40796 14306 40852 14308
rect 40796 14254 40798 14306
rect 40798 14254 40850 14306
rect 40850 14254 40852 14306
rect 40796 14252 40852 14254
rect 41244 14252 41300 14308
rect 41020 12402 41076 12404
rect 41020 12350 41022 12402
rect 41022 12350 41074 12402
rect 41074 12350 41076 12402
rect 41020 12348 41076 12350
rect 40796 11340 40852 11396
rect 39900 9660 39956 9716
rect 39900 9100 39956 9156
rect 40124 8988 40180 9044
rect 40348 8428 40404 8484
rect 40796 7420 40852 7476
rect 41020 9996 41076 10052
rect 41580 12348 41636 12404
rect 41916 14418 41972 14420
rect 41916 14366 41918 14418
rect 41918 14366 41970 14418
rect 41970 14366 41972 14418
rect 41916 14364 41972 14366
rect 42588 14364 42644 14420
rect 42252 14306 42308 14308
rect 42252 14254 42254 14306
rect 42254 14254 42306 14306
rect 42306 14254 42308 14306
rect 42252 14252 42308 14254
rect 41916 14140 41972 14196
rect 42252 12962 42308 12964
rect 42252 12910 42254 12962
rect 42254 12910 42306 12962
rect 42306 12910 42308 12962
rect 42252 12908 42308 12910
rect 41916 11394 41972 11396
rect 41916 11342 41918 11394
rect 41918 11342 41970 11394
rect 41970 11342 41972 11394
rect 41916 11340 41972 11342
rect 42924 16156 42980 16212
rect 43148 16156 43204 16212
rect 42812 15260 42868 15316
rect 42924 15596 42980 15652
rect 43260 15708 43316 15764
rect 43484 15596 43540 15652
rect 43148 15148 43204 15204
rect 43708 15314 43764 15316
rect 43708 15262 43710 15314
rect 43710 15262 43762 15314
rect 43762 15262 43764 15314
rect 43708 15260 43764 15262
rect 43148 12908 43204 12964
rect 43372 15036 43428 15092
rect 43708 15036 43764 15092
rect 43708 12908 43764 12964
rect 42700 10386 42756 10388
rect 42700 10334 42702 10386
rect 42702 10334 42754 10386
rect 42754 10334 42756 10386
rect 42700 10332 42756 10334
rect 41692 10108 41748 10164
rect 41244 9100 41300 9156
rect 41468 8988 41524 9044
rect 41916 9996 41972 10052
rect 42700 9884 42756 9940
rect 42700 9548 42756 9604
rect 44156 20188 44212 20244
rect 44828 16210 44884 16212
rect 44828 16158 44830 16210
rect 44830 16158 44882 16210
rect 44882 16158 44884 16210
rect 44828 16156 44884 16158
rect 44492 15932 44548 15988
rect 43932 15820 43988 15876
rect 44044 15708 44100 15764
rect 44604 15426 44660 15428
rect 44604 15374 44606 15426
rect 44606 15374 44658 15426
rect 44658 15374 44660 15426
rect 44604 15372 44660 15374
rect 44380 15202 44436 15204
rect 44380 15150 44382 15202
rect 44382 15150 44434 15202
rect 44434 15150 44436 15202
rect 44380 15148 44436 15150
rect 44828 11676 44884 11732
rect 44156 10892 44212 10948
rect 43596 9714 43652 9716
rect 43596 9662 43598 9714
rect 43598 9662 43650 9714
rect 43650 9662 43652 9714
rect 43596 9660 43652 9662
rect 41916 9100 41972 9156
rect 42812 8876 42868 8932
rect 42252 8540 42308 8596
rect 41804 7868 41860 7924
rect 42476 7868 42532 7924
rect 41804 6578 41860 6580
rect 41804 6526 41806 6578
rect 41806 6526 41858 6578
rect 41858 6526 41860 6578
rect 41804 6524 41860 6526
rect 42028 6524 42084 6580
rect 37100 4620 37156 4676
rect 36988 4508 37044 4564
rect 33180 4396 33236 4452
rect 33852 4450 33908 4452
rect 33852 4398 33854 4450
rect 33854 4398 33906 4450
rect 33906 4398 33908 4450
rect 33852 4396 33908 4398
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 38892 3724 38948 3780
rect 39788 3724 39844 3780
rect 16156 3276 16212 3332
rect 16940 3330 16996 3332
rect 16940 3278 16942 3330
rect 16942 3278 16994 3330
rect 16994 3278 16996 3330
rect 16940 3276 16996 3278
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 34076 3612 34132 3668
rect 36988 3666 37044 3668
rect 36988 3614 36990 3666
rect 36990 3614 37042 3666
rect 37042 3614 37044 3666
rect 36988 3612 37044 3614
rect 40236 4562 40292 4564
rect 40236 4510 40238 4562
rect 40238 4510 40290 4562
rect 40290 4510 40292 4562
rect 40236 4508 40292 4510
rect 41692 6076 41748 6132
rect 40572 4508 40628 4564
rect 41020 4508 41076 4564
rect 42364 6076 42420 6132
rect 42476 6690 42532 6692
rect 42476 6638 42478 6690
rect 42478 6638 42530 6690
rect 42530 6638 42532 6690
rect 42476 6636 42532 6638
rect 43036 8428 43092 8484
rect 43372 9100 43428 9156
rect 43372 8540 43428 8596
rect 43260 5852 43316 5908
rect 42140 5068 42196 5124
rect 43820 5068 43876 5124
rect 44044 7698 44100 7700
rect 44044 7646 44046 7698
rect 44046 7646 44098 7698
rect 44098 7646 44100 7698
rect 44044 7644 44100 7646
rect 44044 7308 44100 7364
rect 44044 4956 44100 5012
rect 35532 3554 35588 3556
rect 35532 3502 35534 3554
rect 35534 3502 35586 3554
rect 35586 3502 35588 3554
rect 35532 3500 35588 3502
rect 35980 3554 36036 3556
rect 35980 3502 35982 3554
rect 35982 3502 36034 3554
rect 36034 3502 36036 3554
rect 35980 3500 36036 3502
rect 38556 3388 38612 3444
rect 39340 3442 39396 3444
rect 39340 3390 39342 3442
rect 39342 3390 39394 3442
rect 39394 3390 39396 3442
rect 39340 3388 39396 3390
rect 39788 3442 39844 3444
rect 39788 3390 39790 3442
rect 39790 3390 39842 3442
rect 39842 3390 39844 3442
rect 39788 3388 39844 3390
rect 44268 9772 44324 9828
rect 44268 9602 44324 9604
rect 44268 9550 44270 9602
rect 44270 9550 44322 9602
rect 44322 9550 44324 9602
rect 44268 9548 44324 9550
rect 44492 10108 44548 10164
rect 44380 8876 44436 8932
rect 44828 8316 44884 8372
rect 45052 18338 45108 18340
rect 45052 18286 45054 18338
rect 45054 18286 45106 18338
rect 45106 18286 45108 18338
rect 45052 18284 45108 18286
rect 46396 21810 46452 21812
rect 46396 21758 46398 21810
rect 46398 21758 46450 21810
rect 46450 21758 46452 21810
rect 46396 21756 46452 21758
rect 45836 21586 45892 21588
rect 45836 21534 45838 21586
rect 45838 21534 45890 21586
rect 45890 21534 45892 21586
rect 45836 21532 45892 21534
rect 45724 20972 45780 21028
rect 45500 20188 45556 20244
rect 45612 19180 45668 19236
rect 45500 18562 45556 18564
rect 45500 18510 45502 18562
rect 45502 18510 45554 18562
rect 45554 18510 45556 18562
rect 45500 18508 45556 18510
rect 45388 12460 45444 12516
rect 47068 28700 47124 28756
rect 47180 28530 47236 28532
rect 47180 28478 47182 28530
rect 47182 28478 47234 28530
rect 47234 28478 47236 28530
rect 47180 28476 47236 28478
rect 48188 34636 48244 34692
rect 47964 31500 48020 31556
rect 48188 31276 48244 31332
rect 47740 30268 47796 30324
rect 49308 42364 49364 42420
rect 48860 41970 48916 41972
rect 48860 41918 48862 41970
rect 48862 41918 48914 41970
rect 48914 41918 48916 41970
rect 48860 41916 48916 41918
rect 49196 41186 49252 41188
rect 49196 41134 49198 41186
rect 49198 41134 49250 41186
rect 49250 41134 49252 41186
rect 49196 41132 49252 41134
rect 49980 43708 50036 43764
rect 49868 42364 49924 42420
rect 50556 45498 50612 45500
rect 50556 45446 50558 45498
rect 50558 45446 50610 45498
rect 50610 45446 50612 45498
rect 50556 45444 50612 45446
rect 50660 45498 50716 45500
rect 50660 45446 50662 45498
rect 50662 45446 50714 45498
rect 50714 45446 50716 45498
rect 50660 45444 50716 45446
rect 50764 45498 50820 45500
rect 50764 45446 50766 45498
rect 50766 45446 50818 45498
rect 50818 45446 50820 45498
rect 50764 45444 50820 45446
rect 50540 44210 50596 44212
rect 50540 44158 50542 44210
rect 50542 44158 50594 44210
rect 50594 44158 50596 44210
rect 50540 44156 50596 44158
rect 50556 43930 50612 43932
rect 50556 43878 50558 43930
rect 50558 43878 50610 43930
rect 50610 43878 50612 43930
rect 50556 43876 50612 43878
rect 50660 43930 50716 43932
rect 50660 43878 50662 43930
rect 50662 43878 50714 43930
rect 50714 43878 50716 43930
rect 50660 43876 50716 43878
rect 50764 43930 50820 43932
rect 50764 43878 50766 43930
rect 50766 43878 50818 43930
rect 50818 43878 50820 43930
rect 50764 43876 50820 43878
rect 50316 43708 50372 43764
rect 50316 42364 50372 42420
rect 49980 41916 50036 41972
rect 49868 41858 49924 41860
rect 49868 41806 49870 41858
rect 49870 41806 49922 41858
rect 49922 41806 49924 41858
rect 49868 41804 49924 41806
rect 49756 41132 49812 41188
rect 48860 39116 48916 39172
rect 49644 39618 49700 39620
rect 49644 39566 49646 39618
rect 49646 39566 49698 39618
rect 49698 39566 49700 39618
rect 49644 39564 49700 39566
rect 49532 39340 49588 39396
rect 49308 39228 49364 39284
rect 48636 36988 48692 37044
rect 49196 37154 49252 37156
rect 49196 37102 49198 37154
rect 49198 37102 49250 37154
rect 49250 37102 49252 37154
rect 49196 37100 49252 37102
rect 49084 35586 49140 35588
rect 49084 35534 49086 35586
rect 49086 35534 49138 35586
rect 49138 35534 49140 35586
rect 49084 35532 49140 35534
rect 49308 34636 49364 34692
rect 48412 33458 48468 33460
rect 48412 33406 48414 33458
rect 48414 33406 48466 33458
rect 48466 33406 48468 33458
rect 48412 33404 48468 33406
rect 49308 34076 49364 34132
rect 49196 33628 49252 33684
rect 49084 31666 49140 31668
rect 49084 31614 49086 31666
rect 49086 31614 49138 31666
rect 49138 31614 49140 31666
rect 49084 31612 49140 31614
rect 48748 31554 48804 31556
rect 48748 31502 48750 31554
rect 48750 31502 48802 31554
rect 48802 31502 48804 31554
rect 48748 31500 48804 31502
rect 49308 31724 49364 31780
rect 49420 31836 49476 31892
rect 49196 31276 49252 31332
rect 48748 30994 48804 30996
rect 48748 30942 48750 30994
rect 48750 30942 48802 30994
rect 48802 30942 48804 30994
rect 48748 30940 48804 30942
rect 48972 30716 49028 30772
rect 49308 30380 49364 30436
rect 48300 28812 48356 28868
rect 48076 28642 48132 28644
rect 48076 28590 48078 28642
rect 48078 28590 48130 28642
rect 48130 28590 48132 28642
rect 48076 28588 48132 28590
rect 47740 28476 47796 28532
rect 47404 28028 47460 28084
rect 48300 28082 48356 28084
rect 48300 28030 48302 28082
rect 48302 28030 48354 28082
rect 48354 28030 48356 28082
rect 48300 28028 48356 28030
rect 49644 38780 49700 38836
rect 50556 42362 50612 42364
rect 50556 42310 50558 42362
rect 50558 42310 50610 42362
rect 50610 42310 50612 42362
rect 50556 42308 50612 42310
rect 50660 42362 50716 42364
rect 50660 42310 50662 42362
rect 50662 42310 50714 42362
rect 50714 42310 50716 42362
rect 50660 42308 50716 42310
rect 50764 42362 50820 42364
rect 50764 42310 50766 42362
rect 50766 42310 50818 42362
rect 50818 42310 50820 42362
rect 50764 42308 50820 42310
rect 50428 41970 50484 41972
rect 50428 41918 50430 41970
rect 50430 41918 50482 41970
rect 50482 41918 50484 41970
rect 50428 41916 50484 41918
rect 51100 41858 51156 41860
rect 51100 41806 51102 41858
rect 51102 41806 51154 41858
rect 51154 41806 51156 41858
rect 51100 41804 51156 41806
rect 50556 40794 50612 40796
rect 50556 40742 50558 40794
rect 50558 40742 50610 40794
rect 50610 40742 50612 40794
rect 50556 40740 50612 40742
rect 50660 40794 50716 40796
rect 50660 40742 50662 40794
rect 50662 40742 50714 40794
rect 50714 40742 50716 40794
rect 50660 40740 50716 40742
rect 50764 40794 50820 40796
rect 50764 40742 50766 40794
rect 50766 40742 50818 40794
rect 50818 40742 50820 40794
rect 50764 40740 50820 40742
rect 51660 46620 51716 46676
rect 53228 46844 53284 46900
rect 53004 46172 53060 46228
rect 50428 39452 50484 39508
rect 50204 39394 50260 39396
rect 50204 39342 50206 39394
rect 50206 39342 50258 39394
rect 50258 39342 50260 39394
rect 50204 39340 50260 39342
rect 50764 39618 50820 39620
rect 50764 39566 50766 39618
rect 50766 39566 50818 39618
rect 50818 39566 50820 39618
rect 50764 39564 50820 39566
rect 53004 43484 53060 43540
rect 53228 43426 53284 43428
rect 53228 43374 53230 43426
rect 53230 43374 53282 43426
rect 53282 43374 53284 43426
rect 53228 43372 53284 43374
rect 53228 41132 53284 41188
rect 51884 40796 51940 40852
rect 50652 39340 50708 39396
rect 50556 39226 50612 39228
rect 50556 39174 50558 39226
rect 50558 39174 50610 39226
rect 50610 39174 50612 39226
rect 50556 39172 50612 39174
rect 50660 39226 50716 39228
rect 50660 39174 50662 39226
rect 50662 39174 50714 39226
rect 50714 39174 50716 39226
rect 50660 39172 50716 39174
rect 50764 39226 50820 39228
rect 50764 39174 50766 39226
rect 50766 39174 50818 39226
rect 50818 39174 50820 39226
rect 50764 39172 50820 39174
rect 50428 38834 50484 38836
rect 50428 38782 50430 38834
rect 50430 38782 50482 38834
rect 50482 38782 50484 38834
rect 50428 38780 50484 38782
rect 50556 37658 50612 37660
rect 50556 37606 50558 37658
rect 50558 37606 50610 37658
rect 50610 37606 50612 37658
rect 50556 37604 50612 37606
rect 50660 37658 50716 37660
rect 50660 37606 50662 37658
rect 50662 37606 50714 37658
rect 50714 37606 50716 37658
rect 50660 37604 50716 37606
rect 50764 37658 50820 37660
rect 50764 37606 50766 37658
rect 50766 37606 50818 37658
rect 50818 37606 50820 37658
rect 50764 37604 50820 37606
rect 49756 35810 49812 35812
rect 49756 35758 49758 35810
rect 49758 35758 49810 35810
rect 49810 35758 49812 35810
rect 49756 35756 49812 35758
rect 49980 34076 50036 34132
rect 51548 39394 51604 39396
rect 51548 39342 51550 39394
rect 51550 39342 51602 39394
rect 51602 39342 51604 39394
rect 51548 39340 51604 39342
rect 50988 36988 51044 37044
rect 50652 36370 50708 36372
rect 50652 36318 50654 36370
rect 50654 36318 50706 36370
rect 50706 36318 50708 36370
rect 50652 36316 50708 36318
rect 51100 36370 51156 36372
rect 51100 36318 51102 36370
rect 51102 36318 51154 36370
rect 51154 36318 51156 36370
rect 51100 36316 51156 36318
rect 50540 36204 50596 36260
rect 50876 36204 50932 36260
rect 50556 36090 50612 36092
rect 50556 36038 50558 36090
rect 50558 36038 50610 36090
rect 50610 36038 50612 36090
rect 50556 36036 50612 36038
rect 50660 36090 50716 36092
rect 50660 36038 50662 36090
rect 50662 36038 50714 36090
rect 50714 36038 50716 36090
rect 50660 36036 50716 36038
rect 50764 36090 50820 36092
rect 50764 36038 50766 36090
rect 50766 36038 50818 36090
rect 50818 36038 50820 36090
rect 50764 36036 50820 36038
rect 50652 34636 50708 34692
rect 50556 34522 50612 34524
rect 50556 34470 50558 34522
rect 50558 34470 50610 34522
rect 50610 34470 50612 34522
rect 50556 34468 50612 34470
rect 50660 34522 50716 34524
rect 50660 34470 50662 34522
rect 50662 34470 50714 34522
rect 50714 34470 50716 34522
rect 50660 34468 50716 34470
rect 50764 34522 50820 34524
rect 50764 34470 50766 34522
rect 50766 34470 50818 34522
rect 50818 34470 50820 34522
rect 50764 34468 50820 34470
rect 49868 34018 49924 34020
rect 49868 33966 49870 34018
rect 49870 33966 49922 34018
rect 49922 33966 49924 34018
rect 49868 33964 49924 33966
rect 49756 33516 49812 33572
rect 50540 33852 50596 33908
rect 51324 35756 51380 35812
rect 51100 34018 51156 34020
rect 51100 33966 51102 34018
rect 51102 33966 51154 34018
rect 51154 33966 51156 34018
rect 51100 33964 51156 33966
rect 52108 39506 52164 39508
rect 52108 39454 52110 39506
rect 52110 39454 52162 39506
rect 52162 39454 52164 39506
rect 52108 39452 52164 39454
rect 53228 39564 53284 39620
rect 53004 38108 53060 38164
rect 51884 36988 51940 37044
rect 53228 36988 53284 37044
rect 53004 35474 53060 35476
rect 53004 35422 53006 35474
rect 53006 35422 53058 35474
rect 53058 35422 53060 35474
rect 53004 35420 53060 35422
rect 51772 33964 51828 34020
rect 53228 34018 53284 34020
rect 53228 33966 53230 34018
rect 53230 33966 53282 34018
rect 53282 33966 53284 34018
rect 53228 33964 53284 33966
rect 51212 33516 51268 33572
rect 49868 32732 49924 32788
rect 49756 31500 49812 31556
rect 50556 32954 50612 32956
rect 50556 32902 50558 32954
rect 50558 32902 50610 32954
rect 50610 32902 50612 32954
rect 50556 32900 50612 32902
rect 50660 32954 50716 32956
rect 50660 32902 50662 32954
rect 50662 32902 50714 32954
rect 50714 32902 50716 32954
rect 50660 32900 50716 32902
rect 50764 32954 50820 32956
rect 50764 32902 50766 32954
rect 50766 32902 50818 32954
rect 50818 32902 50820 32954
rect 50764 32900 50820 32902
rect 50428 31778 50484 31780
rect 50428 31726 50430 31778
rect 50430 31726 50482 31778
rect 50482 31726 50484 31778
rect 50428 31724 50484 31726
rect 51100 31724 51156 31780
rect 53004 32732 53060 32788
rect 50652 31554 50708 31556
rect 50652 31502 50654 31554
rect 50654 31502 50706 31554
rect 50706 31502 50708 31554
rect 50652 31500 50708 31502
rect 50556 31386 50612 31388
rect 50556 31334 50558 31386
rect 50558 31334 50610 31386
rect 50610 31334 50612 31386
rect 50556 31332 50612 31334
rect 50660 31386 50716 31388
rect 50660 31334 50662 31386
rect 50662 31334 50714 31386
rect 50714 31334 50716 31386
rect 50660 31332 50716 31334
rect 50764 31386 50820 31388
rect 50764 31334 50766 31386
rect 50766 31334 50818 31386
rect 50818 31334 50820 31386
rect 50764 31332 50820 31334
rect 49980 31164 50036 31220
rect 50204 30434 50260 30436
rect 50204 30382 50206 30434
rect 50206 30382 50258 30434
rect 50258 30382 50260 30434
rect 50204 30380 50260 30382
rect 53116 31724 53172 31780
rect 50428 30322 50484 30324
rect 50428 30270 50430 30322
rect 50430 30270 50482 30322
rect 50482 30270 50484 30322
rect 50428 30268 50484 30270
rect 51100 30156 51156 30212
rect 49532 28252 49588 28308
rect 50556 29818 50612 29820
rect 50556 29766 50558 29818
rect 50558 29766 50610 29818
rect 50610 29766 50612 29818
rect 50556 29764 50612 29766
rect 50660 29818 50716 29820
rect 50660 29766 50662 29818
rect 50662 29766 50714 29818
rect 50714 29766 50716 29818
rect 50660 29764 50716 29766
rect 50764 29818 50820 29820
rect 50764 29766 50766 29818
rect 50766 29766 50818 29818
rect 50818 29766 50820 29818
rect 50764 29764 50820 29766
rect 52220 30098 52276 30100
rect 52220 30046 52222 30098
rect 52222 30046 52274 30098
rect 52274 30046 52276 30098
rect 52220 30044 52276 30046
rect 50428 28588 50484 28644
rect 48972 28082 49028 28084
rect 48972 28030 48974 28082
rect 48974 28030 49026 28082
rect 49026 28030 49028 28082
rect 48972 28028 49028 28030
rect 49644 26908 49700 26964
rect 47068 24050 47124 24052
rect 47068 23998 47070 24050
rect 47070 23998 47122 24050
rect 47122 23998 47124 24050
rect 47068 23996 47124 23998
rect 46732 23548 46788 23604
rect 46508 20972 46564 21028
rect 46620 23436 46676 23492
rect 46620 21980 46676 22036
rect 45948 20802 46004 20804
rect 45948 20750 45950 20802
rect 45950 20750 46002 20802
rect 46002 20750 46004 20802
rect 45948 20748 46004 20750
rect 46508 20802 46564 20804
rect 46508 20750 46510 20802
rect 46510 20750 46562 20802
rect 46562 20750 46564 20802
rect 46508 20748 46564 20750
rect 47292 21586 47348 21588
rect 47292 21534 47294 21586
rect 47294 21534 47346 21586
rect 47346 21534 47348 21586
rect 47292 21532 47348 21534
rect 45836 20524 45892 20580
rect 46396 20188 46452 20244
rect 45948 19852 46004 19908
rect 45948 19180 46004 19236
rect 46060 19740 46116 19796
rect 45836 18396 45892 18452
rect 45724 14364 45780 14420
rect 45836 15484 45892 15540
rect 45612 12738 45668 12740
rect 45612 12686 45614 12738
rect 45614 12686 45666 12738
rect 45666 12686 45668 12738
rect 45612 12684 45668 12686
rect 45388 11228 45444 11284
rect 46284 19234 46340 19236
rect 46284 19182 46286 19234
rect 46286 19182 46338 19234
rect 46338 19182 46340 19234
rect 46284 19180 46340 19182
rect 46172 18508 46228 18564
rect 46172 18338 46228 18340
rect 46172 18286 46174 18338
rect 46174 18286 46226 18338
rect 46226 18286 46228 18338
rect 46172 18284 46228 18286
rect 46620 19180 46676 19236
rect 46956 20578 47012 20580
rect 46956 20526 46958 20578
rect 46958 20526 47010 20578
rect 47010 20526 47012 20578
rect 46956 20524 47012 20526
rect 47404 20188 47460 20244
rect 46844 19740 46900 19796
rect 46732 18956 46788 19012
rect 46396 15538 46452 15540
rect 46396 15486 46398 15538
rect 46398 15486 46450 15538
rect 46450 15486 46452 15538
rect 46396 15484 46452 15486
rect 47180 17388 47236 17444
rect 46956 15986 47012 15988
rect 46956 15934 46958 15986
rect 46958 15934 47010 15986
rect 47010 15934 47012 15986
rect 46956 15932 47012 15934
rect 47068 15426 47124 15428
rect 47068 15374 47070 15426
rect 47070 15374 47122 15426
rect 47122 15374 47124 15426
rect 47068 15372 47124 15374
rect 47068 15148 47124 15204
rect 46060 14924 46116 14980
rect 47740 25506 47796 25508
rect 47740 25454 47742 25506
rect 47742 25454 47794 25506
rect 47794 25454 47796 25506
rect 47740 25452 47796 25454
rect 47964 25340 48020 25396
rect 49532 26178 49588 26180
rect 49532 26126 49534 26178
rect 49534 26126 49586 26178
rect 49586 26126 49588 26178
rect 49532 26124 49588 26126
rect 49420 25452 49476 25508
rect 48188 25394 48244 25396
rect 48188 25342 48190 25394
rect 48190 25342 48242 25394
rect 48242 25342 48244 25394
rect 48188 25340 48244 25342
rect 48412 25228 48468 25284
rect 47628 23714 47684 23716
rect 47628 23662 47630 23714
rect 47630 23662 47682 23714
rect 47682 23662 47684 23714
rect 47628 23660 47684 23662
rect 48860 25282 48916 25284
rect 48860 25230 48862 25282
rect 48862 25230 48914 25282
rect 48914 25230 48916 25282
rect 48860 25228 48916 25230
rect 49308 25394 49364 25396
rect 49308 25342 49310 25394
rect 49310 25342 49362 25394
rect 49362 25342 49364 25394
rect 49308 25340 49364 25342
rect 50556 28250 50612 28252
rect 50556 28198 50558 28250
rect 50558 28198 50610 28250
rect 50610 28198 50612 28250
rect 50556 28196 50612 28198
rect 50660 28250 50716 28252
rect 50660 28198 50662 28250
rect 50662 28198 50714 28250
rect 50714 28198 50716 28250
rect 50660 28196 50716 28198
rect 50764 28250 50820 28252
rect 50764 28198 50766 28250
rect 50766 28198 50818 28250
rect 50818 28198 50820 28250
rect 50764 28196 50820 28198
rect 50876 26908 50932 26964
rect 50556 26682 50612 26684
rect 50556 26630 50558 26682
rect 50558 26630 50610 26682
rect 50610 26630 50612 26682
rect 50556 26628 50612 26630
rect 50660 26682 50716 26684
rect 50660 26630 50662 26682
rect 50662 26630 50714 26682
rect 50714 26630 50716 26682
rect 50660 26628 50716 26630
rect 50764 26682 50820 26684
rect 50764 26630 50766 26682
rect 50766 26630 50818 26682
rect 50818 26630 50820 26682
rect 50764 26628 50820 26630
rect 50092 25564 50148 25620
rect 49084 24610 49140 24612
rect 49084 24558 49086 24610
rect 49086 24558 49138 24610
rect 49138 24558 49140 24610
rect 49084 24556 49140 24558
rect 49644 24556 49700 24612
rect 50204 25394 50260 25396
rect 50204 25342 50206 25394
rect 50206 25342 50258 25394
rect 50258 25342 50260 25394
rect 50204 25340 50260 25342
rect 48300 23548 48356 23604
rect 47964 23042 48020 23044
rect 47964 22990 47966 23042
rect 47966 22990 48018 23042
rect 48018 22990 48020 23042
rect 47964 22988 48020 22990
rect 47852 22092 47908 22148
rect 47628 20188 47684 20244
rect 47964 21698 48020 21700
rect 47964 21646 47966 21698
rect 47966 21646 48018 21698
rect 48018 21646 48020 21698
rect 47964 21644 48020 21646
rect 48076 20860 48132 20916
rect 50204 24556 50260 24612
rect 49420 23660 49476 23716
rect 49308 22876 49364 22932
rect 48860 22146 48916 22148
rect 48860 22094 48862 22146
rect 48862 22094 48914 22146
rect 48914 22094 48916 22146
rect 48860 22092 48916 22094
rect 49532 23042 49588 23044
rect 49532 22990 49534 23042
rect 49534 22990 49586 23042
rect 49586 22990 49588 23042
rect 49532 22988 49588 22990
rect 50988 26124 51044 26180
rect 50556 25114 50612 25116
rect 50556 25062 50558 25114
rect 50558 25062 50610 25114
rect 50610 25062 50612 25114
rect 50556 25060 50612 25062
rect 50660 25114 50716 25116
rect 50660 25062 50662 25114
rect 50662 25062 50714 25114
rect 50714 25062 50716 25114
rect 50660 25060 50716 25062
rect 50764 25114 50820 25116
rect 50764 25062 50766 25114
rect 50766 25062 50818 25114
rect 50818 25062 50820 25114
rect 50764 25060 50820 25062
rect 50652 24610 50708 24612
rect 50652 24558 50654 24610
rect 50654 24558 50706 24610
rect 50706 24558 50708 24610
rect 50652 24556 50708 24558
rect 50556 23546 50612 23548
rect 50556 23494 50558 23546
rect 50558 23494 50610 23546
rect 50610 23494 50612 23546
rect 50556 23492 50612 23494
rect 50660 23546 50716 23548
rect 50660 23494 50662 23546
rect 50662 23494 50714 23546
rect 50714 23494 50716 23546
rect 50660 23492 50716 23494
rect 50764 23546 50820 23548
rect 50764 23494 50766 23546
rect 50766 23494 50818 23546
rect 50818 23494 50820 23546
rect 50764 23492 50820 23494
rect 50428 23212 50484 23268
rect 50316 22764 50372 22820
rect 50428 22428 50484 22484
rect 49420 21810 49476 21812
rect 49420 21758 49422 21810
rect 49422 21758 49474 21810
rect 49474 21758 49476 21810
rect 49420 21756 49476 21758
rect 48748 21698 48804 21700
rect 48748 21646 48750 21698
rect 48750 21646 48802 21698
rect 48802 21646 48804 21698
rect 48748 21644 48804 21646
rect 48636 21532 48692 21588
rect 49308 21698 49364 21700
rect 49308 21646 49310 21698
rect 49310 21646 49362 21698
rect 49362 21646 49364 21698
rect 49308 21644 49364 21646
rect 49756 22258 49812 22260
rect 49756 22206 49758 22258
rect 49758 22206 49810 22258
rect 49810 22206 49812 22258
rect 49756 22204 49812 22206
rect 50204 22258 50260 22260
rect 50204 22206 50206 22258
rect 50206 22206 50258 22258
rect 50258 22206 50260 22258
rect 50204 22204 50260 22206
rect 49868 21868 49924 21924
rect 49980 21980 50036 22036
rect 48860 20748 48916 20804
rect 47964 19068 48020 19124
rect 48188 19010 48244 19012
rect 48188 18958 48190 19010
rect 48190 18958 48242 19010
rect 48242 18958 48244 19010
rect 48188 18956 48244 18958
rect 47628 17554 47684 17556
rect 47628 17502 47630 17554
rect 47630 17502 47682 17554
rect 47682 17502 47684 17554
rect 47628 17500 47684 17502
rect 48188 17554 48244 17556
rect 48188 17502 48190 17554
rect 48190 17502 48242 17554
rect 48242 17502 48244 17554
rect 48188 17500 48244 17502
rect 48412 19068 48468 19124
rect 47740 17442 47796 17444
rect 47740 17390 47742 17442
rect 47742 17390 47794 17442
rect 47794 17390 47796 17442
rect 47740 17388 47796 17390
rect 47628 16828 47684 16884
rect 47964 15538 48020 15540
rect 47964 15486 47966 15538
rect 47966 15486 48018 15538
rect 48018 15486 48020 15538
rect 47964 15484 48020 15486
rect 47628 15372 47684 15428
rect 46396 15036 46452 15092
rect 46508 14364 46564 14420
rect 46172 14306 46228 14308
rect 46172 14254 46174 14306
rect 46174 14254 46226 14306
rect 46226 14254 46228 14306
rect 46172 14252 46228 14254
rect 46396 14252 46452 14308
rect 46060 14140 46116 14196
rect 46172 13916 46228 13972
rect 45724 12460 45780 12516
rect 45948 11788 46004 11844
rect 45612 11228 45668 11284
rect 45052 10892 45108 10948
rect 45052 10556 45108 10612
rect 45724 10610 45780 10612
rect 45724 10558 45726 10610
rect 45726 10558 45778 10610
rect 45778 10558 45780 10610
rect 45724 10556 45780 10558
rect 45052 9826 45108 9828
rect 45052 9774 45054 9826
rect 45054 9774 45106 9826
rect 45106 9774 45108 9826
rect 45052 9772 45108 9774
rect 45164 9548 45220 9604
rect 45052 8988 45108 9044
rect 45500 10108 45556 10164
rect 45388 9772 45444 9828
rect 46284 12738 46340 12740
rect 46284 12686 46286 12738
rect 46286 12686 46338 12738
rect 46338 12686 46340 12738
rect 46284 12684 46340 12686
rect 46172 11676 46228 11732
rect 46172 9996 46228 10052
rect 45388 8988 45444 9044
rect 46172 9266 46228 9268
rect 46172 9214 46174 9266
rect 46174 9214 46226 9266
rect 46226 9214 46228 9266
rect 46172 9212 46228 9214
rect 45612 8652 45668 8708
rect 45276 8316 45332 8372
rect 45164 7420 45220 7476
rect 45388 7980 45444 8036
rect 45500 7644 45556 7700
rect 45612 8428 45668 8484
rect 45388 6748 45444 6804
rect 45164 6578 45220 6580
rect 45164 6526 45166 6578
rect 45166 6526 45218 6578
rect 45218 6526 45220 6578
rect 45164 6524 45220 6526
rect 45500 6578 45556 6580
rect 45500 6526 45502 6578
rect 45502 6526 45554 6578
rect 45554 6526 45556 6578
rect 45500 6524 45556 6526
rect 44940 6076 44996 6132
rect 46620 11676 46676 11732
rect 46396 10610 46452 10612
rect 46396 10558 46398 10610
rect 46398 10558 46450 10610
rect 46450 10558 46452 10610
rect 46396 10556 46452 10558
rect 46844 14306 46900 14308
rect 46844 14254 46846 14306
rect 46846 14254 46898 14306
rect 46898 14254 46900 14306
rect 46844 14252 46900 14254
rect 46844 13244 46900 13300
rect 46956 12236 47012 12292
rect 47404 13244 47460 13300
rect 46732 10556 46788 10612
rect 46060 7868 46116 7924
rect 46620 9548 46676 9604
rect 46620 9100 46676 9156
rect 47180 10610 47236 10612
rect 47180 10558 47182 10610
rect 47182 10558 47234 10610
rect 47234 10558 47236 10610
rect 47180 10556 47236 10558
rect 46956 9548 47012 9604
rect 46844 8316 46900 8372
rect 47068 7756 47124 7812
rect 46284 7474 46340 7476
rect 46284 7422 46286 7474
rect 46286 7422 46338 7474
rect 46338 7422 46340 7474
rect 46284 7420 46340 7422
rect 46060 6412 46116 6468
rect 46620 6524 46676 6580
rect 47404 6578 47460 6580
rect 47404 6526 47406 6578
rect 47406 6526 47458 6578
rect 47458 6526 47460 6578
rect 47404 6524 47460 6526
rect 46732 6412 46788 6468
rect 50876 22988 50932 23044
rect 50556 21978 50612 21980
rect 50556 21926 50558 21978
rect 50558 21926 50610 21978
rect 50610 21926 50612 21978
rect 50556 21924 50612 21926
rect 50660 21978 50716 21980
rect 50660 21926 50662 21978
rect 50662 21926 50714 21978
rect 50714 21926 50716 21978
rect 50660 21924 50716 21926
rect 50764 21978 50820 21980
rect 50764 21926 50766 21978
rect 50766 21926 50818 21978
rect 50818 21926 50820 21978
rect 50764 21924 50820 21926
rect 48860 17836 48916 17892
rect 48524 17666 48580 17668
rect 48524 17614 48526 17666
rect 48526 17614 48578 17666
rect 48578 17614 48580 17666
rect 48524 17612 48580 17614
rect 48860 17442 48916 17444
rect 48860 17390 48862 17442
rect 48862 17390 48914 17442
rect 48914 17390 48916 17442
rect 48860 17388 48916 17390
rect 49980 20914 50036 20916
rect 49980 20862 49982 20914
rect 49982 20862 50034 20914
rect 50034 20862 50036 20914
rect 49980 20860 50036 20862
rect 50556 20410 50612 20412
rect 50556 20358 50558 20410
rect 50558 20358 50610 20410
rect 50610 20358 50612 20410
rect 50556 20356 50612 20358
rect 50660 20410 50716 20412
rect 50660 20358 50662 20410
rect 50662 20358 50714 20410
rect 50714 20358 50716 20410
rect 50660 20356 50716 20358
rect 50764 20410 50820 20412
rect 50764 20358 50766 20410
rect 50766 20358 50818 20410
rect 50818 20358 50820 20410
rect 50764 20356 50820 20358
rect 50204 19852 50260 19908
rect 49308 18844 49364 18900
rect 50204 19122 50260 19124
rect 50204 19070 50206 19122
rect 50206 19070 50258 19122
rect 50258 19070 50260 19122
rect 50204 19068 50260 19070
rect 50316 18956 50372 19012
rect 50092 18844 50148 18900
rect 50540 19740 50596 19796
rect 50988 19180 51044 19236
rect 50764 19122 50820 19124
rect 50764 19070 50766 19122
rect 50766 19070 50818 19122
rect 50818 19070 50820 19122
rect 50764 19068 50820 19070
rect 50556 18842 50612 18844
rect 50556 18790 50558 18842
rect 50558 18790 50610 18842
rect 50610 18790 50612 18842
rect 50556 18788 50612 18790
rect 50660 18842 50716 18844
rect 50660 18790 50662 18842
rect 50662 18790 50714 18842
rect 50714 18790 50716 18842
rect 50660 18788 50716 18790
rect 50764 18842 50820 18844
rect 50764 18790 50766 18842
rect 50766 18790 50818 18842
rect 50818 18790 50820 18842
rect 50764 18788 50820 18790
rect 50540 18620 50596 18676
rect 49196 18396 49252 18452
rect 49756 17836 49812 17892
rect 49308 17666 49364 17668
rect 49308 17614 49310 17666
rect 49310 17614 49362 17666
rect 49362 17614 49364 17666
rect 49308 17612 49364 17614
rect 49196 17052 49252 17108
rect 48748 16882 48804 16884
rect 48748 16830 48750 16882
rect 48750 16830 48802 16882
rect 48802 16830 48804 16882
rect 48748 16828 48804 16830
rect 49420 16882 49476 16884
rect 49420 16830 49422 16882
rect 49422 16830 49474 16882
rect 49474 16830 49476 16882
rect 49420 16828 49476 16830
rect 49084 16380 49140 16436
rect 49644 17052 49700 17108
rect 50316 18338 50372 18340
rect 50316 18286 50318 18338
rect 50318 18286 50370 18338
rect 50370 18286 50372 18338
rect 50316 18284 50372 18286
rect 50876 18338 50932 18340
rect 50876 18286 50878 18338
rect 50878 18286 50930 18338
rect 50930 18286 50932 18338
rect 50876 18284 50932 18286
rect 50556 17274 50612 17276
rect 50556 17222 50558 17274
rect 50558 17222 50610 17274
rect 50610 17222 50612 17274
rect 50556 17220 50612 17222
rect 50660 17274 50716 17276
rect 50660 17222 50662 17274
rect 50662 17222 50714 17274
rect 50714 17222 50716 17274
rect 50660 17220 50716 17222
rect 50764 17274 50820 17276
rect 50764 17222 50766 17274
rect 50766 17222 50818 17274
rect 50818 17222 50820 17274
rect 50764 17220 50820 17222
rect 50204 16828 50260 16884
rect 49980 16604 50036 16660
rect 49980 16380 50036 16436
rect 49980 16156 50036 16212
rect 49084 15036 49140 15092
rect 48860 14530 48916 14532
rect 48860 14478 48862 14530
rect 48862 14478 48914 14530
rect 48914 14478 48916 14530
rect 48860 14476 48916 14478
rect 50556 15706 50612 15708
rect 50556 15654 50558 15706
rect 50558 15654 50610 15706
rect 50610 15654 50612 15706
rect 50556 15652 50612 15654
rect 50660 15706 50716 15708
rect 50660 15654 50662 15706
rect 50662 15654 50714 15706
rect 50714 15654 50716 15706
rect 50660 15652 50716 15654
rect 50764 15706 50820 15708
rect 50764 15654 50766 15706
rect 50766 15654 50818 15706
rect 50818 15654 50820 15706
rect 50764 15652 50820 15654
rect 50204 15484 50260 15540
rect 49980 14588 50036 14644
rect 49644 14476 49700 14532
rect 48636 13244 48692 13300
rect 49084 14252 49140 14308
rect 48972 12460 49028 12516
rect 48972 11788 49028 11844
rect 49644 13580 49700 13636
rect 50316 15314 50372 15316
rect 50316 15262 50318 15314
rect 50318 15262 50370 15314
rect 50370 15262 50372 15314
rect 50316 15260 50372 15262
rect 53228 31500 53284 31556
rect 53228 30098 53284 30100
rect 53228 30046 53230 30098
rect 53230 30046 53282 30098
rect 53282 30046 53284 30098
rect 53228 30044 53284 30046
rect 52668 27356 52724 27412
rect 53228 27356 53284 27412
rect 53228 25564 53284 25620
rect 52556 23996 52612 24052
rect 53228 24722 53284 24724
rect 53228 24670 53230 24722
rect 53230 24670 53282 24722
rect 53282 24670 53284 24722
rect 53228 24668 53284 24670
rect 52892 23884 52948 23940
rect 53228 22428 53284 22484
rect 53340 21980 53396 22036
rect 52892 21756 52948 21812
rect 52332 17388 52388 17444
rect 52780 21532 52836 21588
rect 50988 16716 51044 16772
rect 52892 20748 52948 20804
rect 53228 19906 53284 19908
rect 53228 19854 53230 19906
rect 53230 19854 53282 19906
rect 53282 19854 53284 19906
rect 53228 19852 53284 19854
rect 53228 19292 53284 19348
rect 53228 16770 53284 16772
rect 53228 16718 53230 16770
rect 53230 16718 53282 16770
rect 53282 16718 53284 16770
rect 53228 16716 53284 16718
rect 53116 16604 53172 16660
rect 50988 15260 51044 15316
rect 50652 15148 50708 15204
rect 52668 14642 52724 14644
rect 52668 14590 52670 14642
rect 52670 14590 52722 14642
rect 52722 14590 52724 14642
rect 52668 14588 52724 14590
rect 50556 14138 50612 14140
rect 50556 14086 50558 14138
rect 50558 14086 50610 14138
rect 50610 14086 50612 14138
rect 50556 14084 50612 14086
rect 50660 14138 50716 14140
rect 50660 14086 50662 14138
rect 50662 14086 50714 14138
rect 50714 14086 50716 14138
rect 50660 14084 50716 14086
rect 50764 14138 50820 14140
rect 50764 14086 50766 14138
rect 50766 14086 50818 14138
rect 50818 14086 50820 14138
rect 50764 14084 50820 14086
rect 52220 13916 52276 13972
rect 53228 13916 53284 13972
rect 53228 13634 53284 13636
rect 53228 13582 53230 13634
rect 53230 13582 53282 13634
rect 53282 13582 53284 13634
rect 53228 13580 53284 13582
rect 47964 9660 48020 9716
rect 48860 9772 48916 9828
rect 48524 9212 48580 9268
rect 48636 8316 48692 8372
rect 47740 8258 47796 8260
rect 47740 8206 47742 8258
rect 47742 8206 47794 8258
rect 47794 8206 47796 8258
rect 47740 8204 47796 8206
rect 49196 10610 49252 10612
rect 49196 10558 49198 10610
rect 49198 10558 49250 10610
rect 49250 10558 49252 10610
rect 49196 10556 49252 10558
rect 49308 9884 49364 9940
rect 50764 12738 50820 12740
rect 50764 12686 50766 12738
rect 50766 12686 50818 12738
rect 50818 12686 50820 12738
rect 50764 12684 50820 12686
rect 50556 12570 50612 12572
rect 50556 12518 50558 12570
rect 50558 12518 50610 12570
rect 50610 12518 50612 12570
rect 50556 12516 50612 12518
rect 50660 12570 50716 12572
rect 50660 12518 50662 12570
rect 50662 12518 50714 12570
rect 50714 12518 50716 12570
rect 50660 12516 50716 12518
rect 50764 12570 50820 12572
rect 50764 12518 50766 12570
rect 50766 12518 50818 12570
rect 50818 12518 50820 12570
rect 50764 12516 50820 12518
rect 52444 12290 52500 12292
rect 52444 12238 52446 12290
rect 52446 12238 52498 12290
rect 52498 12238 52500 12290
rect 52444 12236 52500 12238
rect 53228 11282 53284 11284
rect 53228 11230 53230 11282
rect 53230 11230 53282 11282
rect 53282 11230 53284 11282
rect 53228 11228 53284 11230
rect 50556 11002 50612 11004
rect 50556 10950 50558 11002
rect 50558 10950 50610 11002
rect 50610 10950 50612 11002
rect 50556 10948 50612 10950
rect 50660 11002 50716 11004
rect 50660 10950 50662 11002
rect 50662 10950 50714 11002
rect 50714 10950 50716 11002
rect 50660 10948 50716 10950
rect 50764 11002 50820 11004
rect 50764 10950 50766 11002
rect 50766 10950 50818 11002
rect 50818 10950 50820 11002
rect 50764 10948 50820 10950
rect 49420 9772 49476 9828
rect 49196 9714 49252 9716
rect 49196 9662 49198 9714
rect 49198 9662 49250 9714
rect 49250 9662 49252 9714
rect 49196 9660 49252 9662
rect 49532 9548 49588 9604
rect 49084 8258 49140 8260
rect 49084 8206 49086 8258
rect 49086 8206 49138 8258
rect 49138 8206 49140 8258
rect 49084 8204 49140 8206
rect 48188 8034 48244 8036
rect 48188 7982 48190 8034
rect 48190 7982 48242 8034
rect 48242 7982 48244 8034
rect 48188 7980 48244 7982
rect 47964 7586 48020 7588
rect 47964 7534 47966 7586
rect 47966 7534 48018 7586
rect 48018 7534 48020 7586
rect 47964 7532 48020 7534
rect 48188 7474 48244 7476
rect 48188 7422 48190 7474
rect 48190 7422 48242 7474
rect 48242 7422 48244 7474
rect 48188 7420 48244 7422
rect 47740 6748 47796 6804
rect 48188 6748 48244 6804
rect 46284 5122 46340 5124
rect 46284 5070 46286 5122
rect 46286 5070 46338 5122
rect 46338 5070 46340 5122
rect 46284 5068 46340 5070
rect 46508 5068 46564 5124
rect 44268 4338 44324 4340
rect 44268 4286 44270 4338
rect 44270 4286 44322 4338
rect 44322 4286 44324 4338
rect 44268 4284 44324 4286
rect 48524 7980 48580 8036
rect 48748 6972 48804 7028
rect 48412 6636 48468 6692
rect 48972 6860 49028 6916
rect 49644 8034 49700 8036
rect 49644 7982 49646 8034
rect 49646 7982 49698 8034
rect 49698 7982 49700 8034
rect 49644 7980 49700 7982
rect 49420 7756 49476 7812
rect 49308 7474 49364 7476
rect 49308 7422 49310 7474
rect 49310 7422 49362 7474
rect 49362 7422 49364 7474
rect 49308 7420 49364 7422
rect 49532 7532 49588 7588
rect 49868 9714 49924 9716
rect 49868 9662 49870 9714
rect 49870 9662 49922 9714
rect 49922 9662 49924 9714
rect 49868 9660 49924 9662
rect 52892 9996 52948 10052
rect 50764 9938 50820 9940
rect 50764 9886 50766 9938
rect 50766 9886 50818 9938
rect 50818 9886 50820 9938
rect 50764 9884 50820 9886
rect 50556 9434 50612 9436
rect 50556 9382 50558 9434
rect 50558 9382 50610 9434
rect 50610 9382 50612 9434
rect 50556 9380 50612 9382
rect 50660 9434 50716 9436
rect 50660 9382 50662 9434
rect 50662 9382 50714 9434
rect 50714 9382 50716 9434
rect 50660 9380 50716 9382
rect 50764 9434 50820 9436
rect 50764 9382 50766 9434
rect 50766 9382 50818 9434
rect 50818 9382 50820 9434
rect 50764 9380 50820 9382
rect 53340 9660 53396 9716
rect 53228 8540 53284 8596
rect 50540 8146 50596 8148
rect 50540 8094 50542 8146
rect 50542 8094 50594 8146
rect 50594 8094 50596 8146
rect 50540 8092 50596 8094
rect 50556 7866 50612 7868
rect 50556 7814 50558 7866
rect 50558 7814 50610 7866
rect 50610 7814 50612 7866
rect 50556 7812 50612 7814
rect 50660 7866 50716 7868
rect 50660 7814 50662 7866
rect 50662 7814 50714 7866
rect 50714 7814 50716 7866
rect 50660 7812 50716 7814
rect 50764 7866 50820 7868
rect 50764 7814 50766 7866
rect 50766 7814 50818 7866
rect 50818 7814 50820 7866
rect 50764 7812 50820 7814
rect 52668 8034 52724 8036
rect 52668 7982 52670 8034
rect 52670 7982 52722 8034
rect 52722 7982 52724 8034
rect 52668 7980 52724 7982
rect 49084 6748 49140 6804
rect 49308 6972 49364 7028
rect 49868 6914 49924 6916
rect 49868 6862 49870 6914
rect 49870 6862 49922 6914
rect 49922 6862 49924 6914
rect 49868 6860 49924 6862
rect 49644 6690 49700 6692
rect 49644 6638 49646 6690
rect 49646 6638 49698 6690
rect 49698 6638 49700 6690
rect 49644 6636 49700 6638
rect 50316 6748 50372 6804
rect 51324 6466 51380 6468
rect 51324 6414 51326 6466
rect 51326 6414 51378 6466
rect 51378 6414 51380 6466
rect 51324 6412 51380 6414
rect 50556 6298 50612 6300
rect 50556 6246 50558 6298
rect 50558 6246 50610 6298
rect 50610 6246 50612 6298
rect 50556 6244 50612 6246
rect 50660 6298 50716 6300
rect 50660 6246 50662 6298
rect 50662 6246 50714 6298
rect 50714 6246 50716 6298
rect 50660 6244 50716 6246
rect 50764 6298 50820 6300
rect 50764 6246 50766 6298
rect 50766 6246 50818 6298
rect 50818 6246 50820 6298
rect 50764 6244 50820 6246
rect 51548 6076 51604 6132
rect 52668 6578 52724 6580
rect 52668 6526 52670 6578
rect 52670 6526 52722 6578
rect 52722 6526 52724 6578
rect 52668 6524 52724 6526
rect 51996 6412 52052 6468
rect 48636 5122 48692 5124
rect 48636 5070 48638 5122
rect 48638 5070 48690 5122
rect 48690 5070 48692 5122
rect 48636 5068 48692 5070
rect 49980 5682 50036 5684
rect 49980 5630 49982 5682
rect 49982 5630 50034 5682
rect 50034 5630 50036 5682
rect 49980 5628 50036 5630
rect 48188 4450 48244 4452
rect 48188 4398 48190 4450
rect 48190 4398 48242 4450
rect 48242 4398 48244 4450
rect 48188 4396 48244 4398
rect 47516 4338 47572 4340
rect 47516 4286 47518 4338
rect 47518 4286 47570 4338
rect 47570 4286 47572 4338
rect 47516 4284 47572 4286
rect 49084 4284 49140 4340
rect 51996 5852 52052 5908
rect 51100 5794 51156 5796
rect 51100 5742 51102 5794
rect 51102 5742 51154 5794
rect 51154 5742 51156 5794
rect 51100 5740 51156 5742
rect 53228 5068 53284 5124
rect 52668 4956 52724 5012
rect 50556 4730 50612 4732
rect 50556 4678 50558 4730
rect 50558 4678 50610 4730
rect 50610 4678 50612 4730
rect 50556 4676 50612 4678
rect 50660 4730 50716 4732
rect 50660 4678 50662 4730
rect 50662 4678 50714 4730
rect 50714 4678 50716 4730
rect 50660 4676 50716 4678
rect 50764 4730 50820 4732
rect 50764 4678 50766 4730
rect 50766 4678 50818 4730
rect 50818 4678 50820 4730
rect 50764 4676 50820 4678
rect 50876 4450 50932 4452
rect 50876 4398 50878 4450
rect 50878 4398 50930 4450
rect 50930 4398 50932 4450
rect 50876 4396 50932 4398
rect 50316 4284 50372 4340
rect 51660 4338 51716 4340
rect 51660 4286 51662 4338
rect 51662 4286 51714 4338
rect 51714 4286 51716 4338
rect 51660 4284 51716 4286
rect 46956 3554 47012 3556
rect 46956 3502 46958 3554
rect 46958 3502 47010 3554
rect 47010 3502 47012 3554
rect 46956 3500 47012 3502
rect 47628 3554 47684 3556
rect 47628 3502 47630 3554
rect 47630 3502 47682 3554
rect 47682 3502 47684 3554
rect 47628 3500 47684 3502
rect 50428 3666 50484 3668
rect 50428 3614 50430 3666
rect 50430 3614 50482 3666
rect 50482 3614 50484 3666
rect 50428 3612 50484 3614
rect 51996 3612 52052 3668
rect 47404 3330 47460 3332
rect 47404 3278 47406 3330
rect 47406 3278 47458 3330
rect 47458 3278 47460 3330
rect 47404 3276 47460 3278
rect 50556 3162 50612 3164
rect 50556 3110 50558 3162
rect 50558 3110 50610 3162
rect 50610 3110 50612 3162
rect 50556 3108 50612 3110
rect 50660 3162 50716 3164
rect 50660 3110 50662 3162
rect 50662 3110 50714 3162
rect 50714 3110 50716 3162
rect 50660 3108 50716 3110
rect 50764 3162 50820 3164
rect 50764 3110 50766 3162
rect 50766 3110 50818 3162
rect 50818 3110 50820 3162
rect 50764 3108 50820 3110
rect 52444 3164 52500 3220
rect 53228 3164 53284 3220
<< metal3 >>
rect 19826 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20110 51772
rect 50546 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50830 51772
rect 54200 51604 55000 51632
rect 51090 51548 51100 51604
rect 51156 51548 55000 51604
rect 54200 51520 55000 51548
rect 49634 51324 49644 51380
rect 49700 51324 50652 51380
rect 50708 51324 51212 51380
rect 51268 51324 51278 51380
rect 50418 51212 50428 51268
rect 50484 51212 51436 51268
rect 51492 51212 51502 51268
rect 4466 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4750 50988
rect 35186 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35470 50988
rect 24556 50540 27692 50596
rect 27748 50540 27758 50596
rect 24556 50484 24612 50540
rect 16370 50428 16380 50484
rect 16436 50428 17724 50484
rect 17780 50428 17790 50484
rect 20738 50428 20748 50484
rect 20804 50428 24108 50484
rect 24164 50428 24174 50484
rect 24546 50428 24556 50484
rect 24612 50428 24622 50484
rect 25106 50428 25116 50484
rect 25172 50428 25900 50484
rect 25956 50428 25966 50484
rect 27346 50428 27356 50484
rect 27412 50428 28588 50484
rect 28644 50428 28654 50484
rect 44146 50428 44156 50484
rect 44212 50428 44940 50484
rect 44996 50428 45006 50484
rect 13682 50316 13692 50372
rect 13748 50316 22764 50372
rect 22820 50316 22830 50372
rect 48738 50316 48748 50372
rect 48804 50316 49980 50372
rect 50036 50316 50046 50372
rect 19826 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20110 50204
rect 50546 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50830 50204
rect 18050 49756 18060 49812
rect 18116 49756 19292 49812
rect 19348 49756 19358 49812
rect 24546 49756 24556 49812
rect 24612 49756 25452 49812
rect 25508 49756 25518 49812
rect 37426 49756 37436 49812
rect 37492 49756 38556 49812
rect 38612 49756 38622 49812
rect 13570 49644 13580 49700
rect 13636 49644 15708 49700
rect 15764 49644 16492 49700
rect 16548 49644 18956 49700
rect 19012 49644 19628 49700
rect 19684 49644 20076 49700
rect 20132 49644 20142 49700
rect 23202 49644 23212 49700
rect 23268 49644 24892 49700
rect 24948 49644 24958 49700
rect 25554 49644 25564 49700
rect 25620 49644 31724 49700
rect 31780 49644 31790 49700
rect 48290 49644 48300 49700
rect 48356 49644 49196 49700
rect 49252 49644 49262 49700
rect 27346 49420 27356 49476
rect 27412 49420 28476 49476
rect 28532 49420 30716 49476
rect 30772 49420 30782 49476
rect 35634 49420 35644 49476
rect 35700 49420 37660 49476
rect 37716 49420 37726 49476
rect 37874 49420 37884 49476
rect 37940 49420 38668 49476
rect 4466 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4750 49420
rect 35186 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35470 49420
rect 27020 49308 27244 49364
rect 27300 49308 27310 49364
rect 35532 49308 38500 49364
rect 27020 49028 27076 49308
rect 35532 49140 35588 49308
rect 32050 49084 32060 49140
rect 32116 49084 35196 49140
rect 35252 49084 35588 49140
rect 38444 49140 38500 49308
rect 38612 49252 38668 49420
rect 38612 49196 41132 49252
rect 41188 49196 41198 49252
rect 50194 49196 50204 49252
rect 50260 49196 50428 49252
rect 50484 49196 50494 49252
rect 38444 49084 38668 49140
rect 38724 49084 39788 49140
rect 39844 49084 39854 49140
rect 50372 49084 53228 49140
rect 53284 49084 53294 49140
rect 50372 49028 50428 49084
rect 19618 48972 19628 49028
rect 19684 48972 25228 49028
rect 25284 48972 26684 49028
rect 26740 48972 26750 49028
rect 27010 48972 27020 49028
rect 27076 48972 27086 49028
rect 38210 48972 38220 49028
rect 38276 48972 38286 49028
rect 38546 48972 38556 49028
rect 38612 48972 40012 49028
rect 40068 48972 40908 49028
rect 40964 48972 40974 49028
rect 48738 48972 48748 49028
rect 48804 48972 49980 49028
rect 50036 48972 50428 49028
rect 38220 48916 38276 48972
rect 54200 48916 55000 48944
rect 18386 48860 18396 48916
rect 18452 48860 19516 48916
rect 19572 48860 20300 48916
rect 20356 48860 20366 48916
rect 36754 48860 36764 48916
rect 36820 48860 37212 48916
rect 37268 48860 37548 48916
rect 37604 48860 37996 48916
rect 38052 48860 38062 48916
rect 38220 48860 38668 48916
rect 38724 48860 41356 48916
rect 41412 48860 41422 48916
rect 47170 48860 47180 48916
rect 47236 48860 48412 48916
rect 48468 48860 48972 48916
rect 49028 48860 49038 48916
rect 51874 48860 51884 48916
rect 51940 48860 55000 48916
rect 54200 48832 55000 48860
rect 19394 48748 19404 48804
rect 19460 48748 20188 48804
rect 20244 48748 20254 48804
rect 27906 48748 27916 48804
rect 27972 48748 29148 48804
rect 29204 48748 30940 48804
rect 30996 48748 33964 48804
rect 34020 48748 35532 48804
rect 35588 48748 36876 48804
rect 36932 48748 36942 48804
rect 38434 48748 38444 48804
rect 38500 48748 39004 48804
rect 39060 48748 40348 48804
rect 40404 48748 40414 48804
rect 46386 48748 46396 48804
rect 46452 48748 46956 48804
rect 47012 48748 48188 48804
rect 48244 48748 48254 48804
rect 32284 48692 32340 48748
rect 24434 48636 24444 48692
rect 24500 48636 25676 48692
rect 25732 48636 27132 48692
rect 27188 48636 31052 48692
rect 31108 48636 31118 48692
rect 32274 48636 32284 48692
rect 32340 48636 32350 48692
rect 19826 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20110 48636
rect 50546 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50830 48636
rect 20626 48524 20636 48580
rect 20692 48524 23436 48580
rect 23492 48524 25004 48580
rect 25060 48524 25070 48580
rect 18498 48412 18508 48468
rect 18564 48412 21532 48468
rect 21588 48412 22204 48468
rect 22260 48412 22270 48468
rect 26562 48412 26572 48468
rect 26628 48412 27132 48468
rect 27188 48412 27198 48468
rect 20402 48300 20412 48356
rect 20468 48300 22092 48356
rect 22148 48300 22158 48356
rect 22306 48300 22316 48356
rect 22372 48300 24332 48356
rect 24388 48300 25564 48356
rect 25620 48300 26908 48356
rect 26964 48300 26974 48356
rect 19394 48188 19404 48244
rect 19460 48188 21644 48244
rect 21700 48188 21710 48244
rect 22642 48188 22652 48244
rect 22708 48188 23100 48244
rect 23156 48188 25228 48244
rect 25284 48188 26236 48244
rect 26292 48188 27580 48244
rect 27636 48188 37996 48244
rect 38052 48188 38062 48244
rect 46834 48188 46844 48244
rect 46900 48188 49308 48244
rect 49364 48188 49980 48244
rect 50036 48188 50046 48244
rect 21410 48076 21420 48132
rect 21476 48076 31612 48132
rect 31668 48076 31678 48132
rect 40114 48076 40124 48132
rect 40180 48076 41020 48132
rect 41076 48076 41804 48132
rect 41860 48076 42476 48132
rect 42532 48076 42542 48132
rect 42914 48076 42924 48132
rect 42980 48076 45500 48132
rect 45556 48076 46172 48132
rect 46228 48076 47180 48132
rect 47236 48076 47246 48132
rect 19282 47964 19292 48020
rect 19348 47964 19740 48020
rect 19796 47964 21308 48020
rect 21364 47964 21374 48020
rect 31938 47964 31948 48020
rect 32004 47964 33180 48020
rect 33236 47964 33246 48020
rect 48178 47964 48188 48020
rect 48244 47964 48972 48020
rect 49028 47964 49038 48020
rect 4466 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4750 47852
rect 35186 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35470 47852
rect 24098 47516 24108 47572
rect 24164 47516 26012 47572
rect 26068 47516 27020 47572
rect 27076 47516 27086 47572
rect 33730 47516 33740 47572
rect 33796 47516 35308 47572
rect 35364 47516 35374 47572
rect 37090 47516 37100 47572
rect 37156 47516 38556 47572
rect 38612 47516 38622 47572
rect 11330 47404 11340 47460
rect 11396 47404 14028 47460
rect 14084 47404 17388 47460
rect 17444 47404 17454 47460
rect 26338 47404 26348 47460
rect 26404 47404 28252 47460
rect 28308 47404 28318 47460
rect 40002 47404 40012 47460
rect 40068 47404 41580 47460
rect 41636 47404 41646 47460
rect 13234 47292 13244 47348
rect 13300 47292 14140 47348
rect 14196 47292 14206 47348
rect 25442 47292 25452 47348
rect 25508 47292 26572 47348
rect 26628 47292 26638 47348
rect 28130 47292 28140 47348
rect 28196 47292 29932 47348
rect 29988 47292 29998 47348
rect 41906 47292 41916 47348
rect 41972 47292 42700 47348
rect 42756 47292 42766 47348
rect 46722 47292 46732 47348
rect 46788 47292 48748 47348
rect 48804 47292 49868 47348
rect 49924 47292 49934 47348
rect 26226 47180 26236 47236
rect 26292 47180 27132 47236
rect 27188 47180 27198 47236
rect 41794 47180 41804 47236
rect 41860 47180 45724 47236
rect 45780 47180 45790 47236
rect 19826 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20110 47068
rect 50546 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50830 47068
rect 15092 46844 21084 46900
rect 21140 46844 21150 46900
rect 27234 46844 27244 46900
rect 27300 46844 27468 46900
rect 27524 46844 30940 46900
rect 30996 46844 32060 46900
rect 32116 46844 32126 46900
rect 48850 46844 48860 46900
rect 48916 46844 53228 46900
rect 53284 46844 53294 46900
rect 15092 46788 15148 46844
rect 12226 46732 12236 46788
rect 12292 46732 14028 46788
rect 14084 46732 15148 46788
rect 20402 46732 20412 46788
rect 20468 46732 20972 46788
rect 21028 46732 21038 46788
rect 23426 46732 23436 46788
rect 23492 46732 23996 46788
rect 24052 46732 24444 46788
rect 24500 46732 24510 46788
rect 26852 46732 33516 46788
rect 33572 46732 33582 46788
rect 26852 46676 26908 46732
rect 12338 46620 12348 46676
rect 12404 46620 13132 46676
rect 13188 46620 13198 46676
rect 19394 46620 19404 46676
rect 19460 46620 20300 46676
rect 20356 46620 26908 46676
rect 28466 46620 28476 46676
rect 28532 46620 30268 46676
rect 30324 46620 30334 46676
rect 38332 46620 38892 46676
rect 38948 46620 40012 46676
rect 40068 46620 40078 46676
rect 42466 46620 42476 46676
rect 42532 46620 47068 46676
rect 47124 46620 48188 46676
rect 48244 46620 48748 46676
rect 48804 46620 48814 46676
rect 50372 46620 50988 46676
rect 51044 46620 51660 46676
rect 51716 46620 51726 46676
rect 38332 46564 38388 46620
rect 50372 46564 50428 46620
rect 12786 46508 12796 46564
rect 12852 46508 13356 46564
rect 13412 46508 13422 46564
rect 22530 46508 22540 46564
rect 22596 46508 29932 46564
rect 29988 46508 29998 46564
rect 36194 46508 36204 46564
rect 36260 46508 37100 46564
rect 37156 46508 37166 46564
rect 38322 46508 38332 46564
rect 38388 46508 38398 46564
rect 38612 46508 38780 46564
rect 38836 46508 38846 46564
rect 44146 46508 44156 46564
rect 44212 46508 46508 46564
rect 46564 46508 46574 46564
rect 49298 46508 49308 46564
rect 49364 46508 50428 46564
rect 38612 46452 38668 46508
rect 37538 46396 37548 46452
rect 37604 46396 38668 46452
rect 42242 46396 42252 46452
rect 42308 46396 42924 46452
rect 42980 46396 44380 46452
rect 44436 46396 44446 46452
rect 4466 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4750 46284
rect 35186 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35470 46284
rect 54200 46228 55000 46256
rect 18722 46172 18732 46228
rect 18788 46172 19180 46228
rect 19236 46172 19246 46228
rect 52994 46172 53004 46228
rect 53060 46172 55000 46228
rect 54200 46144 55000 46172
rect 13122 45948 13132 46004
rect 13188 45948 14252 46004
rect 14308 45948 14318 46004
rect 14018 45836 14028 45892
rect 14084 45836 14588 45892
rect 14644 45836 14654 45892
rect 22418 45836 22428 45892
rect 22484 45836 23436 45892
rect 23492 45836 23502 45892
rect 38210 45836 38220 45892
rect 38276 45836 40236 45892
rect 40292 45836 40302 45892
rect 40562 45836 40572 45892
rect 40628 45836 41132 45892
rect 41188 45836 42028 45892
rect 42084 45836 43260 45892
rect 43316 45836 43326 45892
rect 49298 45836 49308 45892
rect 49364 45836 50204 45892
rect 50260 45836 50270 45892
rect 40236 45780 40292 45836
rect 36978 45724 36988 45780
rect 37044 45724 37884 45780
rect 37940 45724 37950 45780
rect 38658 45724 38668 45780
rect 38724 45724 39564 45780
rect 39620 45724 39630 45780
rect 40236 45724 41468 45780
rect 41524 45724 42364 45780
rect 42420 45724 42980 45780
rect 43138 45724 43148 45780
rect 43204 45724 43820 45780
rect 43876 45724 43886 45780
rect 42924 45668 42980 45724
rect 12450 45612 12460 45668
rect 12516 45612 14252 45668
rect 14308 45612 14318 45668
rect 15922 45612 15932 45668
rect 15988 45612 16492 45668
rect 16548 45612 19180 45668
rect 19236 45612 19246 45668
rect 24658 45612 24668 45668
rect 24724 45612 25452 45668
rect 25508 45612 25518 45668
rect 36306 45612 36316 45668
rect 36372 45612 39788 45668
rect 39844 45612 40236 45668
rect 40292 45612 40302 45668
rect 42914 45612 42924 45668
rect 42980 45612 42990 45668
rect 49186 45612 49196 45668
rect 49252 45612 49868 45668
rect 49924 45612 49934 45668
rect 11554 45500 11564 45556
rect 11620 45500 12348 45556
rect 12404 45500 12414 45556
rect 13906 45500 13916 45556
rect 13972 45500 15148 45556
rect 15204 45500 16380 45556
rect 16436 45500 16940 45556
rect 16996 45500 17006 45556
rect 22642 45500 22652 45556
rect 22708 45500 24780 45556
rect 24836 45500 24846 45556
rect 42690 45500 42700 45556
rect 42756 45500 43148 45556
rect 43204 45500 44044 45556
rect 44100 45500 44110 45556
rect 19826 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20110 45500
rect 50546 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50830 45500
rect 12226 45388 12236 45444
rect 12292 45388 13580 45444
rect 13636 45388 16268 45444
rect 16324 45388 16334 45444
rect 21970 45388 21980 45444
rect 22036 45388 22876 45444
rect 22932 45388 23772 45444
rect 23828 45388 23838 45444
rect 30146 45388 30156 45444
rect 30212 45388 30940 45444
rect 30996 45388 31006 45444
rect 9426 45276 9436 45332
rect 9492 45276 11564 45332
rect 11620 45276 11630 45332
rect 18610 45276 18620 45332
rect 18676 45276 19628 45332
rect 19684 45276 19694 45332
rect 23202 45276 23212 45332
rect 23268 45276 25228 45332
rect 25284 45276 25294 45332
rect 32274 45276 32284 45332
rect 32340 45276 37324 45332
rect 37380 45276 38780 45332
rect 38836 45276 38846 45332
rect 42242 45276 42252 45332
rect 42308 45276 43372 45332
rect 43428 45276 46060 45332
rect 46116 45276 46620 45332
rect 46676 45276 46686 45332
rect 19068 45220 19124 45276
rect 11778 45164 11788 45220
rect 11844 45164 12124 45220
rect 12180 45164 12190 45220
rect 18050 45164 18060 45220
rect 18116 45164 18844 45220
rect 18900 45164 18910 45220
rect 19058 45164 19068 45220
rect 19124 45164 19162 45220
rect 34850 45164 34860 45220
rect 34916 45164 38332 45220
rect 38388 45164 38892 45220
rect 38948 45164 38958 45220
rect 39442 45164 39452 45220
rect 39508 45164 48748 45220
rect 48804 45164 50092 45220
rect 50148 45164 50158 45220
rect 14130 45052 14140 45108
rect 14196 45052 18284 45108
rect 18340 45052 21868 45108
rect 21924 45052 21934 45108
rect 34626 45052 34636 45108
rect 34692 45052 35756 45108
rect 35812 45052 35822 45108
rect 37426 45052 37436 45108
rect 37492 45052 38444 45108
rect 38500 45052 38510 45108
rect 40002 45052 40012 45108
rect 40068 45052 40908 45108
rect 40964 45052 40974 45108
rect 48290 45052 48300 45108
rect 48356 45052 48972 45108
rect 49028 45052 49038 45108
rect 15362 44940 15372 44996
rect 15428 44940 23996 44996
rect 24052 44940 24556 44996
rect 24612 44940 24622 44996
rect 28354 44940 28364 44996
rect 28420 44940 31500 44996
rect 31556 44940 31566 44996
rect 32834 44940 32844 44996
rect 32900 44940 35420 44996
rect 35476 44940 35486 44996
rect 43250 44940 43260 44996
rect 43316 44940 44492 44996
rect 44548 44940 44558 44996
rect 19058 44828 19068 44884
rect 19124 44828 19852 44884
rect 19908 44828 19918 44884
rect 23426 44828 23436 44884
rect 23492 44828 33292 44884
rect 33348 44828 33358 44884
rect 34290 44828 34300 44884
rect 34356 44828 34366 44884
rect 34300 44772 34356 44828
rect 24658 44716 24668 44772
rect 24724 44716 34356 44772
rect 4466 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4750 44716
rect 35186 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35470 44716
rect 18274 44604 18284 44660
rect 18340 44604 19740 44660
rect 19796 44604 28364 44660
rect 28420 44604 28430 44660
rect 49074 44604 49084 44660
rect 49140 44604 49756 44660
rect 49812 44604 49822 44660
rect 16594 44492 16604 44548
rect 16660 44492 17276 44548
rect 17332 44492 17342 44548
rect 17714 44380 17724 44436
rect 17780 44380 18396 44436
rect 18452 44380 18620 44436
rect 18676 44380 18686 44436
rect 32050 44380 32060 44436
rect 32116 44380 32844 44436
rect 32900 44380 32910 44436
rect 33394 44380 33404 44436
rect 33460 44380 33964 44436
rect 34020 44380 34860 44436
rect 34916 44380 34926 44436
rect 16146 44268 16156 44324
rect 16212 44268 16828 44324
rect 16884 44268 18172 44324
rect 18228 44268 18238 44324
rect 25218 44268 25228 44324
rect 25284 44268 25564 44324
rect 25620 44268 25630 44324
rect 34178 44268 34188 44324
rect 34244 44268 35756 44324
rect 35812 44268 35822 44324
rect 14466 44156 14476 44212
rect 14532 44156 18396 44212
rect 18452 44156 22540 44212
rect 22596 44156 23492 44212
rect 49634 44156 49644 44212
rect 49700 44156 50540 44212
rect 50596 44156 50606 44212
rect 23436 44100 23492 44156
rect 19506 44044 19516 44100
rect 19572 44044 20300 44100
rect 20356 44044 20366 44100
rect 22082 44044 22092 44100
rect 22148 44044 23212 44100
rect 23268 44044 23278 44100
rect 23426 44044 23436 44100
rect 23492 44044 23502 44100
rect 26226 44044 26236 44100
rect 26292 44044 27020 44100
rect 27076 44044 27086 44100
rect 38658 44044 38668 44100
rect 38724 44044 39564 44100
rect 39620 44044 39630 44100
rect 19826 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20110 43932
rect 50546 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50830 43932
rect 18722 43708 18732 43764
rect 18788 43708 19292 43764
rect 19348 43708 19358 43764
rect 21410 43708 21420 43764
rect 21476 43708 25116 43764
rect 25172 43708 27468 43764
rect 27524 43708 27534 43764
rect 33730 43708 33740 43764
rect 33796 43708 34188 43764
rect 34244 43708 34254 43764
rect 49970 43708 49980 43764
rect 50036 43708 50316 43764
rect 50372 43708 50382 43764
rect 11778 43596 11788 43652
rect 11844 43596 14028 43652
rect 14084 43596 14094 43652
rect 14252 43596 20748 43652
rect 20804 43596 20814 43652
rect 10882 43484 10892 43540
rect 10948 43484 11452 43540
rect 11508 43484 12516 43540
rect 12460 43428 12516 43484
rect 14252 43428 14308 43596
rect 54200 43540 55000 43568
rect 18946 43484 18956 43540
rect 19012 43484 20412 43540
rect 20468 43484 20478 43540
rect 25890 43484 25900 43540
rect 25956 43484 27132 43540
rect 27188 43484 27198 43540
rect 28578 43484 28588 43540
rect 28644 43484 29260 43540
rect 29316 43484 29326 43540
rect 33954 43484 33964 43540
rect 34020 43484 47516 43540
rect 47572 43484 47582 43540
rect 52994 43484 53004 43540
rect 53060 43484 55000 43540
rect 54200 43456 55000 43484
rect 9650 43372 9660 43428
rect 9716 43372 12012 43428
rect 12068 43372 12078 43428
rect 12460 43372 14308 43428
rect 17042 43372 17052 43428
rect 17108 43372 18508 43428
rect 18564 43372 18574 43428
rect 27234 43372 27244 43428
rect 27300 43372 29708 43428
rect 29764 43372 29774 43428
rect 34066 43372 34076 43428
rect 34132 43372 34860 43428
rect 34916 43372 34926 43428
rect 47170 43372 47180 43428
rect 47236 43372 48300 43428
rect 48356 43372 48972 43428
rect 49028 43372 49038 43428
rect 49186 43372 49196 43428
rect 49252 43372 53228 43428
rect 53284 43372 53294 43428
rect 12674 43260 12684 43316
rect 12740 43260 26012 43316
rect 26068 43260 27356 43316
rect 27412 43260 28588 43316
rect 28644 43260 28654 43316
rect 29362 43260 29372 43316
rect 29428 43260 36988 43316
rect 37044 43260 37054 43316
rect 4466 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4750 43148
rect 35186 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35470 43148
rect 14018 43036 14028 43092
rect 14084 43036 14588 43092
rect 14644 43036 14812 43092
rect 14868 43036 14878 43092
rect 36418 42924 36428 42980
rect 36484 42924 38332 42980
rect 38388 42924 38668 42980
rect 38724 42924 48748 42980
rect 48804 42924 48814 42980
rect 12226 42812 12236 42868
rect 12292 42812 13020 42868
rect 13076 42812 13086 42868
rect 41346 42812 41356 42868
rect 41412 42812 43148 42868
rect 43204 42812 43214 42868
rect 43922 42812 43932 42868
rect 43988 42812 44828 42868
rect 44884 42812 45388 42868
rect 45444 42812 45948 42868
rect 46004 42812 46014 42868
rect 36978 42700 36988 42756
rect 37044 42700 37772 42756
rect 37828 42700 38780 42756
rect 38836 42700 39340 42756
rect 39396 42700 39406 42756
rect 40338 42700 40348 42756
rect 40404 42700 43820 42756
rect 43876 42700 44268 42756
rect 44324 42700 46956 42756
rect 47012 42700 47022 42756
rect 12562 42588 12572 42644
rect 12628 42588 13804 42644
rect 13860 42588 13870 42644
rect 14466 42588 14476 42644
rect 14532 42588 14924 42644
rect 14980 42588 14990 42644
rect 38994 42588 39004 42644
rect 39060 42588 39676 42644
rect 39732 42588 39900 42644
rect 39956 42588 43484 42644
rect 43540 42588 43550 42644
rect 15092 42308 15148 42532
rect 15204 42476 15214 42532
rect 32722 42476 32732 42532
rect 32788 42476 33292 42532
rect 33348 42476 34076 42532
rect 34132 42476 34142 42532
rect 30034 42364 30044 42420
rect 30100 42364 30492 42420
rect 30548 42364 49308 42420
rect 49364 42364 49868 42420
rect 49924 42364 50316 42420
rect 50372 42364 50382 42420
rect 19826 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20110 42364
rect 50546 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50830 42364
rect 14802 42252 14812 42308
rect 14868 42252 15148 42308
rect 14130 42140 14140 42196
rect 14196 42140 15036 42196
rect 15092 42140 15102 42196
rect 33170 42140 33180 42196
rect 33236 42140 38444 42196
rect 38500 42140 38510 42196
rect 14578 42028 14588 42084
rect 14644 42028 15148 42084
rect 15204 42028 15214 42084
rect 23212 42028 23884 42084
rect 23940 42028 23950 42084
rect 23212 41972 23268 42028
rect 16370 41916 16380 41972
rect 16436 41916 22988 41972
rect 23044 41916 23268 41972
rect 23426 41916 23436 41972
rect 23492 41916 23772 41972
rect 23828 41916 26124 41972
rect 26180 41916 26190 41972
rect 46946 41916 46956 41972
rect 47012 41916 48076 41972
rect 48132 41916 48860 41972
rect 48916 41916 49980 41972
rect 50036 41916 50428 41972
rect 50484 41916 50494 41972
rect 5058 41804 5068 41860
rect 5124 41804 8316 41860
rect 8372 41804 8876 41860
rect 8932 41804 9884 41860
rect 9940 41804 9950 41860
rect 23436 41804 24668 41860
rect 24724 41804 27356 41860
rect 27412 41804 31948 41860
rect 32004 41804 32014 41860
rect 44258 41804 44268 41860
rect 44324 41804 44940 41860
rect 44996 41804 45276 41860
rect 45332 41804 45342 41860
rect 49858 41804 49868 41860
rect 49924 41804 51100 41860
rect 51156 41804 51166 41860
rect 23436 41748 23492 41804
rect 23426 41692 23436 41748
rect 23492 41692 23502 41748
rect 32172 41692 33292 41748
rect 33348 41692 33358 41748
rect 32172 41636 32228 41692
rect 19506 41580 19516 41636
rect 19572 41580 32172 41636
rect 32228 41580 32238 41636
rect 4466 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4750 41580
rect 35186 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35470 41580
rect 23986 41468 23996 41524
rect 24052 41468 26348 41524
rect 26404 41468 26414 41524
rect 18050 41356 18060 41412
rect 18116 41356 26796 41412
rect 26852 41356 26862 41412
rect 22978 41244 22988 41300
rect 23044 41244 24220 41300
rect 24276 41244 24286 41300
rect 26002 41244 26012 41300
rect 26068 41244 27916 41300
rect 27972 41244 27982 41300
rect 29138 41244 29148 41300
rect 29204 41244 32396 41300
rect 32452 41244 33516 41300
rect 33572 41244 35756 41300
rect 35812 41244 36652 41300
rect 36708 41244 36718 41300
rect 14690 41132 14700 41188
rect 14756 41132 15372 41188
rect 15428 41132 15438 41188
rect 23650 41132 23660 41188
rect 23716 41132 26572 41188
rect 26628 41132 26638 41188
rect 49186 41132 49196 41188
rect 49252 41132 49756 41188
rect 49812 41132 53228 41188
rect 53284 41132 53294 41188
rect 34290 41020 34300 41076
rect 34356 41020 37100 41076
rect 37156 41020 37166 41076
rect 40226 41020 40236 41076
rect 40292 41020 41132 41076
rect 41188 41020 41198 41076
rect 44258 41020 44268 41076
rect 44324 41020 45836 41076
rect 45892 41020 45902 41076
rect 15138 40908 15148 40964
rect 15204 40908 15596 40964
rect 15652 40908 15662 40964
rect 22418 40908 22428 40964
rect 22484 40908 23996 40964
rect 24052 40908 24062 40964
rect 45714 40908 45724 40964
rect 45780 40908 47404 40964
rect 47460 40908 47470 40964
rect 54200 40852 55000 40880
rect 51874 40796 51884 40852
rect 51940 40796 55000 40852
rect 19826 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20110 40796
rect 50546 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50830 40796
rect 54200 40768 55000 40796
rect 22082 40684 22092 40740
rect 22148 40684 22652 40740
rect 22708 40684 23436 40740
rect 23492 40684 28588 40740
rect 28644 40684 28654 40740
rect 22306 40572 22316 40628
rect 22372 40572 23324 40628
rect 23380 40572 23390 40628
rect 38882 40572 38892 40628
rect 38948 40572 40012 40628
rect 40068 40572 42028 40628
rect 42084 40572 42094 40628
rect 19730 40460 19740 40516
rect 19796 40460 25452 40516
rect 25508 40460 25518 40516
rect 35298 40460 35308 40516
rect 35364 40460 38108 40516
rect 38164 40460 43708 40516
rect 43764 40460 44492 40516
rect 44548 40460 44558 40516
rect 16706 40348 16716 40404
rect 16772 40348 18620 40404
rect 18676 40348 19068 40404
rect 19124 40348 19628 40404
rect 19684 40348 19694 40404
rect 23314 40348 23324 40404
rect 23380 40348 24556 40404
rect 24612 40348 24622 40404
rect 25890 40348 25900 40404
rect 25956 40348 29148 40404
rect 29204 40348 29214 40404
rect 39974 40348 40012 40404
rect 40068 40348 40078 40404
rect 40226 40348 40236 40404
rect 40292 40348 40796 40404
rect 40852 40348 40862 40404
rect 12450 40236 12460 40292
rect 12516 40236 15260 40292
rect 15316 40236 15326 40292
rect 20850 40236 20860 40292
rect 20916 40236 21868 40292
rect 21924 40236 21934 40292
rect 32162 40236 32172 40292
rect 32228 40236 33292 40292
rect 33348 40236 38332 40292
rect 38388 40236 38398 40292
rect 42354 40236 42364 40292
rect 42420 40236 43932 40292
rect 43988 40236 43998 40292
rect 4466 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4750 40012
rect 35186 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35470 40012
rect 8418 39788 8428 39844
rect 8484 39788 9548 39844
rect 9604 39788 9614 39844
rect 41458 39788 41468 39844
rect 41524 39788 43036 39844
rect 43092 39788 43102 39844
rect 5030 39676 5068 39732
rect 5124 39676 5134 39732
rect 9762 39676 9772 39732
rect 9828 39676 12796 39732
rect 12852 39676 15148 39732
rect 15204 39676 15214 39732
rect 15474 39676 15484 39732
rect 15540 39676 16380 39732
rect 16436 39676 16446 39732
rect 38434 39676 38444 39732
rect 38500 39676 39900 39732
rect 39956 39676 39966 39732
rect 9314 39564 9324 39620
rect 9380 39564 10220 39620
rect 10276 39564 10286 39620
rect 13570 39564 13580 39620
rect 13636 39564 16716 39620
rect 16772 39564 16782 39620
rect 36418 39564 36428 39620
rect 36484 39564 37100 39620
rect 37156 39564 38668 39620
rect 40338 39564 40348 39620
rect 40404 39564 41356 39620
rect 41412 39564 45612 39620
rect 45668 39564 45678 39620
rect 46274 39564 46284 39620
rect 46340 39564 46844 39620
rect 46900 39564 49644 39620
rect 49700 39564 49710 39620
rect 50754 39564 50764 39620
rect 50820 39564 53228 39620
rect 53284 39564 53294 39620
rect 4946 39452 4956 39508
rect 5012 39452 6524 39508
rect 6580 39452 8092 39508
rect 8148 39452 8158 39508
rect 9426 39452 9436 39508
rect 9492 39452 10668 39508
rect 10724 39452 10734 39508
rect 38612 39396 38668 39564
rect 44258 39452 44268 39508
rect 44324 39452 46060 39508
rect 46116 39452 46126 39508
rect 50418 39452 50428 39508
rect 50484 39452 52108 39508
rect 52164 39452 52174 39508
rect 51548 39396 51604 39452
rect 5058 39340 5068 39396
rect 5124 39340 5516 39396
rect 5572 39340 5582 39396
rect 6066 39340 6076 39396
rect 6132 39340 7196 39396
rect 7252 39340 8316 39396
rect 8372 39340 8382 39396
rect 38612 39340 39228 39396
rect 39284 39340 39294 39396
rect 40898 39340 40908 39396
rect 40964 39340 45276 39396
rect 45332 39340 45342 39396
rect 49522 39340 49532 39396
rect 49588 39340 50204 39396
rect 50260 39340 50270 39396
rect 50372 39340 50652 39396
rect 50708 39340 50718 39396
rect 51538 39340 51548 39396
rect 51604 39340 51614 39396
rect 6300 39284 6356 39340
rect 50372 39284 50428 39340
rect 6290 39228 6300 39284
rect 6356 39228 6366 39284
rect 9874 39228 9884 39284
rect 9940 39228 11004 39284
rect 11060 39228 11070 39284
rect 36194 39228 36204 39284
rect 36260 39228 37212 39284
rect 37268 39228 38556 39284
rect 38612 39228 38622 39284
rect 49298 39228 49308 39284
rect 49364 39228 50428 39284
rect 19826 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20110 39228
rect 50546 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50830 39228
rect 46946 39116 46956 39172
rect 47012 39116 48860 39172
rect 48916 39116 48926 39172
rect 7970 39004 7980 39060
rect 8036 39004 8316 39060
rect 8372 39004 9772 39060
rect 9828 39004 9838 39060
rect 43026 39004 43036 39060
rect 43092 39004 46396 39060
rect 46452 39004 47292 39060
rect 47348 39004 47358 39060
rect 18162 38892 18172 38948
rect 18228 38892 19740 38948
rect 19796 38892 19806 38948
rect 9734 38780 9772 38836
rect 9828 38780 9838 38836
rect 16594 38780 16604 38836
rect 16660 38780 17612 38836
rect 17668 38780 17678 38836
rect 45714 38780 45724 38836
rect 45780 38780 46284 38836
rect 46340 38780 46350 38836
rect 49634 38780 49644 38836
rect 49700 38780 50428 38836
rect 50484 38780 50494 38836
rect 42802 38668 42812 38724
rect 42868 38668 43932 38724
rect 43988 38668 43998 38724
rect 5394 38556 5404 38612
rect 5460 38556 6412 38612
rect 6468 38556 8988 38612
rect 9044 38556 9054 38612
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 16818 38332 16828 38388
rect 16884 38332 19068 38388
rect 19124 38332 19134 38388
rect 5852 38220 6300 38276
rect 6356 38220 6366 38276
rect 5852 38164 5908 38220
rect 54200 38164 55000 38192
rect 5842 38108 5852 38164
rect 5908 38108 5918 38164
rect 52994 38108 53004 38164
rect 53060 38108 55000 38164
rect 54200 38080 55000 38108
rect 6038 37996 6076 38052
rect 6132 37996 6142 38052
rect 15922 37996 15932 38052
rect 15988 37996 18060 38052
rect 18116 37996 18126 38052
rect 24434 37996 24444 38052
rect 24500 37996 25788 38052
rect 25844 37996 25854 38052
rect 26338 37996 26348 38052
rect 26404 37996 26908 38052
rect 26964 37996 26974 38052
rect 37538 37996 37548 38052
rect 37604 37996 40908 38052
rect 40964 37996 40974 38052
rect 5954 37884 5964 37940
rect 6020 37884 7196 37940
rect 7252 37884 7262 37940
rect 17714 37884 17724 37940
rect 17780 37884 20636 37940
rect 20692 37884 20702 37940
rect 28578 37884 28588 37940
rect 28644 37884 29484 37940
rect 29540 37884 29550 37940
rect 34290 37884 34300 37940
rect 34356 37884 37100 37940
rect 37156 37884 37166 37940
rect 5058 37772 5068 37828
rect 5124 37772 6076 37828
rect 6132 37772 6142 37828
rect 9874 37772 9884 37828
rect 9940 37772 10444 37828
rect 10500 37772 10510 37828
rect 28466 37772 28476 37828
rect 28532 37772 29260 37828
rect 29316 37772 29326 37828
rect 8866 37660 8876 37716
rect 8932 37660 9548 37716
rect 9604 37660 9772 37716
rect 9828 37660 9838 37716
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 50546 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50830 37660
rect 7858 37548 7868 37604
rect 7924 37548 10780 37604
rect 10836 37548 10846 37604
rect 26450 37548 26460 37604
rect 26516 37548 28084 37604
rect 5506 37436 5516 37492
rect 5572 37436 6412 37492
rect 6468 37436 7420 37492
rect 7476 37436 7486 37492
rect 28028 37380 28084 37548
rect 29362 37436 29372 37492
rect 29428 37436 31948 37492
rect 32004 37436 32014 37492
rect 25330 37324 25340 37380
rect 25396 37324 26796 37380
rect 26852 37324 26862 37380
rect 28018 37324 28028 37380
rect 28084 37324 28094 37380
rect 42354 37324 42364 37380
rect 42420 37324 44044 37380
rect 44100 37324 44110 37380
rect 6066 37212 6076 37268
rect 6132 37212 8764 37268
rect 8820 37212 9324 37268
rect 9380 37212 9390 37268
rect 10210 37212 10220 37268
rect 10276 37212 11788 37268
rect 11844 37212 11854 37268
rect 19030 37212 19068 37268
rect 19124 37212 19134 37268
rect 26226 37212 26236 37268
rect 26292 37212 28924 37268
rect 28980 37212 28990 37268
rect 2482 37100 2492 37156
rect 2548 37100 5068 37156
rect 5124 37100 5134 37156
rect 6514 37100 6524 37156
rect 6580 37100 8316 37156
rect 8372 37100 8382 37156
rect 10994 37100 11004 37156
rect 11060 37100 13468 37156
rect 13524 37100 14364 37156
rect 14420 37100 14430 37156
rect 33730 37100 33740 37156
rect 33796 37100 36428 37156
rect 36484 37100 37100 37156
rect 37156 37100 37548 37156
rect 37604 37100 37614 37156
rect 38770 37100 38780 37156
rect 38836 37100 40348 37156
rect 40404 37100 40414 37156
rect 46946 37100 46956 37156
rect 47012 37100 49196 37156
rect 49252 37100 49262 37156
rect 4610 36988 4620 37044
rect 4676 36988 6972 37044
rect 7028 36988 7038 37044
rect 9650 36988 9660 37044
rect 9716 36988 13916 37044
rect 13972 36988 16268 37044
rect 16324 36988 16334 37044
rect 39778 36988 39788 37044
rect 39844 36988 42028 37044
rect 42084 36988 48188 37044
rect 48244 36988 48636 37044
rect 48692 36988 48702 37044
rect 50978 36988 50988 37044
rect 51044 36988 51884 37044
rect 51940 36988 53228 37044
rect 53284 36988 53294 37044
rect 22866 36876 22876 36932
rect 22932 36876 26908 36932
rect 26964 36876 26974 36932
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 5954 36652 5964 36708
rect 6020 36652 6076 36708
rect 6132 36652 6142 36708
rect 38994 36652 39004 36708
rect 39060 36652 39676 36708
rect 39732 36652 39742 36708
rect 18274 36540 18284 36596
rect 18340 36540 18732 36596
rect 18788 36540 18798 36596
rect 38210 36540 38220 36596
rect 38276 36540 38892 36596
rect 38948 36540 38958 36596
rect 8306 36428 8316 36484
rect 8372 36428 9436 36484
rect 9492 36428 9502 36484
rect 12898 36428 12908 36484
rect 12964 36428 17724 36484
rect 17780 36428 17790 36484
rect 19142 36428 19180 36484
rect 19236 36428 19246 36484
rect 20626 36428 20636 36484
rect 20692 36428 21644 36484
rect 21700 36428 21710 36484
rect 45266 36428 45276 36484
rect 45332 36428 46172 36484
rect 46228 36428 46238 36484
rect 6066 36316 6076 36372
rect 6132 36316 9100 36372
rect 9156 36316 9166 36372
rect 15474 36316 15484 36372
rect 15540 36316 16044 36372
rect 16100 36316 20076 36372
rect 20132 36316 21868 36372
rect 21924 36316 22316 36372
rect 22372 36316 24668 36372
rect 24724 36316 36204 36372
rect 36260 36316 37324 36372
rect 37380 36316 37390 36372
rect 44034 36316 44044 36372
rect 44100 36316 46060 36372
rect 46116 36316 46126 36372
rect 50642 36316 50652 36372
rect 50708 36316 51100 36372
rect 51156 36316 51166 36372
rect 28466 36204 28476 36260
rect 28532 36204 29148 36260
rect 29204 36204 29214 36260
rect 39330 36204 39340 36260
rect 39396 36204 39788 36260
rect 39844 36204 40012 36260
rect 40068 36204 40078 36260
rect 50530 36204 50540 36260
rect 50596 36204 50876 36260
rect 50932 36204 50942 36260
rect 28130 36092 28140 36148
rect 28196 36092 40460 36148
rect 40516 36092 40526 36148
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 50546 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50830 36092
rect 26852 35980 39340 36036
rect 39396 35980 39406 36036
rect 26852 35924 26908 35980
rect 1810 35868 1820 35924
rect 1876 35868 4844 35924
rect 4900 35868 5068 35924
rect 5124 35868 5134 35924
rect 10882 35868 10892 35924
rect 10948 35868 11676 35924
rect 11732 35868 26908 35924
rect 35746 35868 35756 35924
rect 35812 35868 38892 35924
rect 38948 35868 38958 35924
rect 43474 35756 43484 35812
rect 43540 35756 44492 35812
rect 44548 35756 44558 35812
rect 49746 35756 49756 35812
rect 49812 35756 51324 35812
rect 51380 35756 51390 35812
rect 38210 35644 38220 35700
rect 38276 35644 46284 35700
rect 46340 35644 46350 35700
rect 16594 35532 16604 35588
rect 16660 35532 19292 35588
rect 19348 35532 20748 35588
rect 20804 35532 20814 35588
rect 40898 35532 40908 35588
rect 40964 35532 47068 35588
rect 47124 35532 49084 35588
rect 49140 35532 49150 35588
rect 54200 35476 55000 35504
rect 52994 35420 53004 35476
rect 53060 35420 55000 35476
rect 54200 35392 55000 35420
rect 30258 35308 30268 35364
rect 30324 35308 32732 35364
rect 32788 35308 33068 35364
rect 33124 35308 33516 35364
rect 33572 35308 33582 35364
rect 40226 35308 40236 35364
rect 40292 35308 45948 35364
rect 46004 35308 46014 35364
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 30268 35252 30324 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 8530 35196 8540 35252
rect 8596 35196 18508 35252
rect 18564 35196 18574 35252
rect 28690 35196 28700 35252
rect 28756 35196 29260 35252
rect 29316 35196 30324 35252
rect 5058 35084 5068 35140
rect 5124 35084 5404 35140
rect 5460 35084 5470 35140
rect 29138 34972 29148 35028
rect 29204 34972 32172 35028
rect 32228 34972 35756 35028
rect 35812 34972 35822 35028
rect 36530 34972 36540 35028
rect 36596 34972 39340 35028
rect 39396 34972 42812 35028
rect 42868 34972 43932 35028
rect 43988 34972 44828 35028
rect 44884 34972 44894 35028
rect 6962 34860 6972 34916
rect 7028 34860 9548 34916
rect 9604 34860 14364 34916
rect 14420 34860 14430 34916
rect 14802 34860 14812 34916
rect 14868 34860 15148 34916
rect 20626 34860 20636 34916
rect 20692 34860 22204 34916
rect 22260 34860 24556 34916
rect 24612 34860 24622 34916
rect 28354 34860 28364 34916
rect 28420 34860 36204 34916
rect 36260 34860 38332 34916
rect 38388 34860 38398 34916
rect 40786 34860 40796 34916
rect 40852 34860 41468 34916
rect 41524 34860 41534 34916
rect 2482 34748 2492 34804
rect 2548 34748 5740 34804
rect 5796 34748 5806 34804
rect 15092 34692 15148 34860
rect 15092 34636 15484 34692
rect 15540 34636 16604 34692
rect 16660 34636 16670 34692
rect 18834 34636 18844 34692
rect 18900 34636 19404 34692
rect 19460 34636 20188 34692
rect 20244 34636 24220 34692
rect 24276 34636 24286 34692
rect 24882 34636 24892 34692
rect 24948 34636 25452 34692
rect 25508 34636 25518 34692
rect 28364 34580 28420 34860
rect 35970 34636 35980 34692
rect 36036 34636 37100 34692
rect 37156 34636 37166 34692
rect 41906 34636 41916 34692
rect 41972 34636 43148 34692
rect 43204 34636 47404 34692
rect 47460 34636 47470 34692
rect 48178 34636 48188 34692
rect 48244 34636 49308 34692
rect 49364 34636 50652 34692
rect 50708 34636 50718 34692
rect 5058 34524 5068 34580
rect 5124 34524 5236 34580
rect 24658 34524 24668 34580
rect 24724 34524 28420 34580
rect 5180 34132 5236 34524
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 50546 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50830 34524
rect 36978 34412 36988 34468
rect 37044 34412 37884 34468
rect 37940 34412 37950 34468
rect 7186 34300 7196 34356
rect 7252 34300 8092 34356
rect 8148 34300 8876 34356
rect 8932 34300 8942 34356
rect 33170 34300 33180 34356
rect 33236 34300 33852 34356
rect 33908 34300 33918 34356
rect 38612 34300 45500 34356
rect 45556 34300 45566 34356
rect 18722 34188 18732 34244
rect 18788 34188 27132 34244
rect 27188 34188 30380 34244
rect 30436 34188 30446 34244
rect 5170 34076 5180 34132
rect 5236 34076 5246 34132
rect 10546 34076 10556 34132
rect 10612 34076 11116 34132
rect 11172 34076 13804 34132
rect 13860 34076 13870 34132
rect 23762 34076 23772 34132
rect 23828 34076 24836 34132
rect 24780 34020 24836 34076
rect 38612 34020 38668 34300
rect 38882 34076 38892 34132
rect 38948 34076 39900 34132
rect 39956 34076 42140 34132
rect 42196 34076 42700 34132
rect 42756 34076 43708 34132
rect 43764 34076 43774 34132
rect 49298 34076 49308 34132
rect 49364 34076 49980 34132
rect 50036 34076 50046 34132
rect 17938 33964 17948 34020
rect 18004 33964 19180 34020
rect 19236 33964 19246 34020
rect 20738 33964 20748 34020
rect 20804 33964 23324 34020
rect 23380 33964 23996 34020
rect 24052 33964 24062 34020
rect 24770 33964 24780 34020
rect 24836 33964 26012 34020
rect 26068 33964 38668 34020
rect 49858 33964 49868 34020
rect 49924 33964 51100 34020
rect 51156 33964 51166 34020
rect 51762 33964 51772 34020
rect 51828 33964 53228 34020
rect 53284 33964 53294 34020
rect 51772 33908 51828 33964
rect 30370 33852 30380 33908
rect 30436 33852 30940 33908
rect 30996 33852 33068 33908
rect 33124 33852 35868 33908
rect 35924 33852 35934 33908
rect 50530 33852 50540 33908
rect 50596 33852 51828 33908
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 20514 33628 20524 33684
rect 20580 33628 20692 33684
rect 45938 33628 45948 33684
rect 46004 33628 49196 33684
rect 49252 33628 49262 33684
rect 15092 33516 15484 33572
rect 15540 33516 15550 33572
rect 18946 33516 18956 33572
rect 19012 33516 20412 33572
rect 20468 33516 20478 33572
rect 5730 33292 5740 33348
rect 5796 33292 6412 33348
rect 6468 33292 6478 33348
rect 15026 33292 15036 33348
rect 15092 33292 15148 33516
rect 20636 33460 20692 33628
rect 42466 33516 42476 33572
rect 42532 33516 43372 33572
rect 43428 33516 43438 33572
rect 49746 33516 49756 33572
rect 49812 33516 51212 33572
rect 51268 33516 51278 33572
rect 19618 33404 19628 33460
rect 19684 33404 20692 33460
rect 41010 33404 41020 33460
rect 41076 33404 41468 33460
rect 41524 33404 41534 33460
rect 41794 33404 41804 33460
rect 41860 33404 48412 33460
rect 48468 33404 48478 33460
rect 19394 33292 19404 33348
rect 19460 33292 19964 33348
rect 20020 33292 21532 33348
rect 21588 33292 26908 33348
rect 29698 33292 29708 33348
rect 29764 33292 30268 33348
rect 30324 33292 33180 33348
rect 33236 33292 33852 33348
rect 33908 33292 33918 33348
rect 39442 33292 39452 33348
rect 39508 33292 45612 33348
rect 45668 33292 45678 33348
rect 26852 33236 26908 33292
rect 9874 33180 9884 33236
rect 9940 33180 10668 33236
rect 10724 33180 10734 33236
rect 21634 33180 21644 33236
rect 21700 33180 22764 33236
rect 22820 33180 22830 33236
rect 26852 33180 33740 33236
rect 33796 33180 34300 33236
rect 34356 33180 35756 33236
rect 35812 33180 35822 33236
rect 5954 33068 5964 33124
rect 6020 33068 6636 33124
rect 6692 33068 6702 33124
rect 9426 33068 9436 33124
rect 9492 33068 10220 33124
rect 10276 33068 10286 33124
rect 10444 33068 20860 33124
rect 20916 33068 20926 33124
rect 23426 33068 23436 33124
rect 23492 33068 24108 33124
rect 24164 33068 24174 33124
rect 29138 33068 29148 33124
rect 29204 33068 29596 33124
rect 29652 33068 29662 33124
rect 30482 33068 30492 33124
rect 30548 33068 31276 33124
rect 31332 33068 32844 33124
rect 32900 33068 32910 33124
rect 10444 33012 10500 33068
rect 8306 32956 8316 33012
rect 8372 32956 8764 33012
rect 8820 32956 10500 33012
rect 15026 32956 15036 33012
rect 15092 32956 15372 33012
rect 15428 32956 15438 33012
rect 20290 32956 20300 33012
rect 20356 32956 41804 33012
rect 41860 32956 41870 33012
rect 43362 32956 43372 33012
rect 43428 32956 43932 33012
rect 43988 32956 43998 33012
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 50546 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50830 32956
rect 4610 32844 4620 32900
rect 4676 32844 6412 32900
rect 6468 32844 6478 32900
rect 8866 32844 8876 32900
rect 8932 32844 18284 32900
rect 18340 32844 18844 32900
rect 18900 32844 18910 32900
rect 54200 32788 55000 32816
rect 6738 32732 6748 32788
rect 6804 32732 8316 32788
rect 8372 32732 8382 32788
rect 16594 32732 16604 32788
rect 16660 32732 25452 32788
rect 25508 32732 26236 32788
rect 26292 32732 26302 32788
rect 43586 32732 43596 32788
rect 43652 32732 49868 32788
rect 49924 32732 49934 32788
rect 52994 32732 53004 32788
rect 53060 32732 55000 32788
rect 54200 32704 55000 32732
rect 5282 32620 5292 32676
rect 5348 32620 6076 32676
rect 6132 32620 6142 32676
rect 16146 32620 16156 32676
rect 16212 32620 19068 32676
rect 19124 32620 19134 32676
rect 24098 32620 24108 32676
rect 24164 32620 30380 32676
rect 30436 32620 31500 32676
rect 31556 32620 31566 32676
rect 39890 32620 39900 32676
rect 39956 32620 40460 32676
rect 40516 32620 40526 32676
rect 5842 32508 5852 32564
rect 5908 32508 7084 32564
rect 7140 32508 7980 32564
rect 8036 32508 8046 32564
rect 14354 32508 14364 32564
rect 14420 32508 14812 32564
rect 14868 32508 14878 32564
rect 19506 32508 19516 32564
rect 19572 32508 19852 32564
rect 19908 32508 19918 32564
rect 22978 32508 22988 32564
rect 23044 32508 23548 32564
rect 23604 32508 26908 32564
rect 30482 32508 30492 32564
rect 30548 32508 30828 32564
rect 30884 32508 32284 32564
rect 32340 32508 32350 32564
rect 33170 32508 33180 32564
rect 33236 32508 33516 32564
rect 33572 32508 35308 32564
rect 35364 32508 38780 32564
rect 38836 32508 38846 32564
rect 26852 32452 26908 32508
rect 2482 32396 2492 32452
rect 2548 32396 5404 32452
rect 5460 32396 5470 32452
rect 8530 32396 8540 32452
rect 8596 32396 13020 32452
rect 13076 32396 13692 32452
rect 13748 32396 13758 32452
rect 16930 32396 16940 32452
rect 16996 32396 17724 32452
rect 17780 32396 17790 32452
rect 26852 32396 30940 32452
rect 30996 32396 31948 32452
rect 32004 32396 32014 32452
rect 34402 32396 34412 32452
rect 34468 32396 35980 32452
rect 36036 32396 36046 32452
rect 39442 32396 39452 32452
rect 39508 32396 45612 32452
rect 45668 32396 45678 32452
rect 21634 32284 21644 32340
rect 21700 32284 32788 32340
rect 35522 32284 35532 32340
rect 35588 32284 42588 32340
rect 42644 32284 43148 32340
rect 43204 32284 43214 32340
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 25330 32060 25340 32116
rect 25396 32060 29260 32116
rect 29316 32060 29326 32116
rect 32732 32004 32788 32284
rect 37426 32172 37436 32228
rect 37492 32172 42924 32228
rect 42980 32172 42990 32228
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 33730 32060 33740 32116
rect 33796 32060 34300 32116
rect 34356 32060 34366 32116
rect 43586 32060 43596 32116
rect 43652 32060 45164 32116
rect 45220 32060 45230 32116
rect 10546 31948 10556 32004
rect 10612 31948 13356 32004
rect 13412 31948 13422 32004
rect 25442 31948 25452 32004
rect 25508 31948 25518 32004
rect 26226 31948 26236 32004
rect 26292 31948 28364 32004
rect 28420 31948 28430 32004
rect 29894 31948 29932 32004
rect 29988 31948 29998 32004
rect 32732 31948 40236 32004
rect 40292 31948 40908 32004
rect 40964 31948 40974 32004
rect 25452 31892 25508 31948
rect 1698 31836 1708 31892
rect 1764 31836 4844 31892
rect 4900 31836 11116 31892
rect 11172 31836 11182 31892
rect 14578 31836 14588 31892
rect 14644 31836 15148 31892
rect 16594 31836 16604 31892
rect 16660 31836 18508 31892
rect 18564 31836 18574 31892
rect 23426 31836 23436 31892
rect 23492 31836 25508 31892
rect 28140 31836 33516 31892
rect 33572 31836 33582 31892
rect 34738 31836 34748 31892
rect 34804 31836 35084 31892
rect 35140 31836 35150 31892
rect 49410 31836 49420 31892
rect 49476 31836 51156 31892
rect 15092 31780 15148 31836
rect 28140 31780 28196 31836
rect 51100 31780 51156 31836
rect 6514 31724 6524 31780
rect 6580 31724 7532 31780
rect 7588 31724 9100 31780
rect 9156 31724 9166 31780
rect 15092 31724 28196 31780
rect 28354 31724 28364 31780
rect 28420 31724 32508 31780
rect 32564 31724 37100 31780
rect 37156 31724 37166 31780
rect 39666 31724 39676 31780
rect 39732 31724 39900 31780
rect 39956 31724 40348 31780
rect 40404 31724 41020 31780
rect 41076 31724 41086 31780
rect 42802 31724 42812 31780
rect 42868 31724 43372 31780
rect 43428 31724 43708 31780
rect 43764 31724 43774 31780
rect 44146 31724 44156 31780
rect 44212 31724 49308 31780
rect 49364 31724 49374 31780
rect 50372 31668 50428 31780
rect 50484 31724 50494 31780
rect 51090 31724 51100 31780
rect 51156 31724 53116 31780
rect 53172 31724 53182 31780
rect 5954 31612 5964 31668
rect 6020 31612 6748 31668
rect 6804 31612 8652 31668
rect 8708 31612 8718 31668
rect 23650 31612 23660 31668
rect 23716 31612 25788 31668
rect 25844 31612 25854 31668
rect 28242 31612 28252 31668
rect 28308 31612 42252 31668
rect 42308 31612 42700 31668
rect 42756 31612 42766 31668
rect 49074 31612 49084 31668
rect 49140 31612 50428 31668
rect 5618 31500 5628 31556
rect 5684 31500 6188 31556
rect 6244 31500 6254 31556
rect 9314 31500 9324 31556
rect 9380 31500 9884 31556
rect 9940 31500 9950 31556
rect 13570 31500 13580 31556
rect 13636 31500 17836 31556
rect 17892 31500 20300 31556
rect 20356 31500 25452 31556
rect 25508 31500 25518 31556
rect 31938 31500 31948 31556
rect 32004 31500 32396 31556
rect 32452 31500 33292 31556
rect 33348 31500 33358 31556
rect 33506 31500 33516 31556
rect 33572 31500 34636 31556
rect 34692 31500 35196 31556
rect 35252 31500 38108 31556
rect 38164 31500 38174 31556
rect 44370 31500 44380 31556
rect 44436 31500 45164 31556
rect 45220 31500 47964 31556
rect 48020 31500 48748 31556
rect 48804 31500 48814 31556
rect 49746 31500 49756 31556
rect 49812 31500 50652 31556
rect 50708 31500 53228 31556
rect 53284 31500 53294 31556
rect 6290 31388 6300 31444
rect 6356 31388 6412 31444
rect 6468 31388 6860 31444
rect 6916 31388 6926 31444
rect 24322 31388 24332 31444
rect 24388 31388 42812 31444
rect 42868 31388 42878 31444
rect 43362 31388 43372 31444
rect 43428 31388 43820 31444
rect 43876 31388 43886 31444
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 50546 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50830 31388
rect 24434 31276 24444 31332
rect 24500 31276 25004 31332
rect 25060 31276 25070 31332
rect 33842 31276 33852 31332
rect 33908 31276 34748 31332
rect 34804 31276 34814 31332
rect 37090 31276 37100 31332
rect 37156 31276 37548 31332
rect 37604 31276 37614 31332
rect 48178 31276 48188 31332
rect 48244 31276 49196 31332
rect 49252 31276 49262 31332
rect 36978 31164 36988 31220
rect 37044 31164 37054 31220
rect 43810 31164 43820 31220
rect 43876 31164 49980 31220
rect 50036 31164 50046 31220
rect 36988 31108 37044 31164
rect 9202 31052 9212 31108
rect 9268 31052 10108 31108
rect 10164 31052 10556 31108
rect 10612 31052 10622 31108
rect 24210 31052 24220 31108
rect 24276 31052 24556 31108
rect 24612 31052 25116 31108
rect 25172 31052 37772 31108
rect 37828 31052 37838 31108
rect 43698 31052 43708 31108
rect 43764 31052 44044 31108
rect 44100 31052 44828 31108
rect 44884 31052 44894 31108
rect 6962 30940 6972 30996
rect 7028 30940 8092 30996
rect 8148 30940 8876 30996
rect 8932 30940 8942 30996
rect 14130 30940 14140 30996
rect 14196 30940 17948 30996
rect 18004 30940 18014 30996
rect 18498 30940 18508 30996
rect 18564 30940 24668 30996
rect 24724 30940 25228 30996
rect 25284 30940 25294 30996
rect 37874 30940 37884 30996
rect 37940 30940 39116 30996
rect 39172 30940 39182 30996
rect 43026 30940 43036 30996
rect 43092 30940 43102 30996
rect 45154 30940 45164 30996
rect 45220 30940 48748 30996
rect 48804 30940 48814 30996
rect 43036 30884 43092 30940
rect 5618 30828 5628 30884
rect 5684 30828 6412 30884
rect 6468 30828 6478 30884
rect 16146 30828 16156 30884
rect 16212 30828 16716 30884
rect 16772 30828 21980 30884
rect 22036 30828 22046 30884
rect 25778 30828 25788 30884
rect 25844 30828 26460 30884
rect 26516 30828 33740 30884
rect 33796 30828 33806 30884
rect 34962 30828 34972 30884
rect 35028 30828 35196 30884
rect 35252 30828 36204 30884
rect 36260 30828 36270 30884
rect 36530 30828 36540 30884
rect 36596 30828 43092 30884
rect 7074 30716 7084 30772
rect 7140 30716 15596 30772
rect 15652 30716 15662 30772
rect 39218 30716 39228 30772
rect 39284 30716 48972 30772
rect 49028 30716 49038 30772
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 30146 30492 30156 30548
rect 30212 30492 30716 30548
rect 30772 30492 30782 30548
rect 8642 30380 8652 30436
rect 8708 30380 9548 30436
rect 9604 30380 9614 30436
rect 23874 30380 23884 30436
rect 23940 30380 35532 30436
rect 35588 30380 35598 30436
rect 49298 30380 49308 30436
rect 49364 30380 50204 30436
rect 50260 30380 50270 30436
rect 9762 30268 9772 30324
rect 9828 30268 10220 30324
rect 10276 30268 10668 30324
rect 10724 30268 13468 30324
rect 13524 30268 13534 30324
rect 33282 30268 33292 30324
rect 33348 30268 38220 30324
rect 38276 30268 38286 30324
rect 38994 30268 39004 30324
rect 39060 30268 40908 30324
rect 40964 30268 47740 30324
rect 47796 30268 47806 30324
rect 50418 30268 50428 30324
rect 50484 30268 51156 30324
rect 51100 30212 51156 30268
rect 13346 30156 13356 30212
rect 13412 30156 17724 30212
rect 17780 30156 17790 30212
rect 20290 30156 20300 30212
rect 20356 30156 21868 30212
rect 21924 30156 21934 30212
rect 25554 30156 25564 30212
rect 25620 30156 26236 30212
rect 26292 30156 26302 30212
rect 26852 30156 29372 30212
rect 29428 30156 29820 30212
rect 29876 30156 32396 30212
rect 32452 30156 32462 30212
rect 34626 30156 34636 30212
rect 34692 30156 35532 30212
rect 35588 30156 35598 30212
rect 42578 30156 42588 30212
rect 42644 30156 47068 30212
rect 47124 30156 47292 30212
rect 47348 30156 47358 30212
rect 51090 30156 51100 30212
rect 51156 30156 51166 30212
rect 18162 30044 18172 30100
rect 18228 30044 20636 30100
rect 20692 30044 22540 30100
rect 22596 30044 23324 30100
rect 23380 30044 23390 30100
rect 4946 29932 4956 29988
rect 5012 29932 10108 29988
rect 10164 29932 10174 29988
rect 20402 29932 20412 29988
rect 20468 29932 21420 29988
rect 21476 29932 21486 29988
rect 23762 29932 23772 29988
rect 23828 29932 24556 29988
rect 24612 29932 24622 29988
rect 26852 29876 26908 30156
rect 54200 30100 55000 30128
rect 31154 30044 31164 30100
rect 31220 30044 31836 30100
rect 31892 30044 31902 30100
rect 37986 30044 37996 30100
rect 38052 30044 39452 30100
rect 39508 30044 47068 30100
rect 47124 30044 47134 30100
rect 52210 30044 52220 30100
rect 52276 30044 53228 30100
rect 53284 30044 55000 30100
rect 54200 30016 55000 30044
rect 30706 29932 30716 29988
rect 30772 29932 31500 29988
rect 31556 29932 33628 29988
rect 33684 29932 33694 29988
rect 33954 29932 33964 29988
rect 34020 29932 34412 29988
rect 34468 29932 35084 29988
rect 35140 29932 41132 29988
rect 41188 29932 42028 29988
rect 42084 29932 42094 29988
rect 22418 29820 22428 29876
rect 22484 29820 25340 29876
rect 25396 29820 26908 29876
rect 27346 29820 27356 29876
rect 27412 29820 35756 29876
rect 35812 29820 36428 29876
rect 36484 29820 36494 29876
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 50546 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50830 29820
rect 36978 29708 36988 29764
rect 37044 29708 42028 29764
rect 42084 29708 42588 29764
rect 42644 29708 42654 29764
rect 5282 29596 5292 29652
rect 5348 29596 7308 29652
rect 7364 29596 14812 29652
rect 14868 29596 14878 29652
rect 23202 29596 23212 29652
rect 23268 29596 25228 29652
rect 25284 29596 25294 29652
rect 33730 29596 33740 29652
rect 33796 29596 37884 29652
rect 37940 29596 38444 29652
rect 38500 29596 38510 29652
rect 38994 29596 39004 29652
rect 39060 29596 44940 29652
rect 44996 29596 45006 29652
rect 6066 29484 6076 29540
rect 6132 29484 8204 29540
rect 8260 29484 8270 29540
rect 20290 29484 20300 29540
rect 20356 29484 22876 29540
rect 22932 29484 22942 29540
rect 39638 29484 39676 29540
rect 39732 29484 39742 29540
rect 40338 29484 40348 29540
rect 40404 29484 41244 29540
rect 41300 29484 42140 29540
rect 42196 29484 42206 29540
rect 7308 29316 7364 29484
rect 17490 29372 17500 29428
rect 17556 29372 18844 29428
rect 18900 29372 18910 29428
rect 32386 29372 32396 29428
rect 32452 29372 36316 29428
rect 36372 29372 36382 29428
rect 38994 29372 39004 29428
rect 39060 29372 40684 29428
rect 40740 29372 40750 29428
rect 39564 29316 39620 29372
rect 2818 29260 2828 29316
rect 2884 29260 5292 29316
rect 5348 29260 5358 29316
rect 7298 29260 7308 29316
rect 7364 29260 7374 29316
rect 15092 29260 16828 29316
rect 16884 29260 16894 29316
rect 17826 29260 17836 29316
rect 17892 29260 26124 29316
rect 26180 29260 26460 29316
rect 26516 29260 26526 29316
rect 39554 29260 39564 29316
rect 39620 29260 39630 29316
rect 15092 29204 15148 29260
rect 4610 29148 4620 29204
rect 4676 29148 6860 29204
rect 6916 29148 15148 29204
rect 15362 29148 15372 29204
rect 15428 29148 15932 29204
rect 15988 29148 28924 29204
rect 28980 29148 28990 29204
rect 38210 29148 38220 29204
rect 38276 29148 39340 29204
rect 39396 29148 39406 29204
rect 20402 29036 20412 29092
rect 20468 29036 21420 29092
rect 21476 29036 31164 29092
rect 31220 29036 31230 29092
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 15092 28924 25116 28980
rect 25172 28924 26180 28980
rect 26450 28924 26460 28980
rect 26516 28924 30380 28980
rect 30436 28924 30446 28980
rect 4722 28812 4732 28868
rect 4788 28812 5740 28868
rect 5796 28812 5806 28868
rect 15092 28644 15148 28924
rect 26124 28868 26180 28924
rect 19590 28812 19628 28868
rect 19684 28812 19694 28868
rect 26124 28812 28140 28868
rect 28196 28812 28206 28868
rect 28354 28812 28364 28868
rect 28420 28812 29372 28868
rect 29428 28812 29438 28868
rect 32162 28812 32172 28868
rect 32228 28812 37548 28868
rect 37604 28812 37614 28868
rect 38994 28812 39004 28868
rect 39060 28812 41972 28868
rect 42914 28812 42924 28868
rect 42980 28812 48300 28868
rect 48356 28812 48366 28868
rect 32172 28756 32228 28812
rect 41916 28756 41972 28812
rect 19170 28700 19180 28756
rect 19236 28700 19740 28756
rect 19796 28700 21756 28756
rect 21812 28700 21822 28756
rect 25778 28700 25788 28756
rect 25844 28700 26236 28756
rect 26292 28700 26908 28756
rect 26964 28700 27356 28756
rect 27412 28700 27422 28756
rect 29596 28700 32228 28756
rect 36194 28700 36204 28756
rect 36260 28700 37660 28756
rect 37716 28700 41132 28756
rect 41188 28700 41198 28756
rect 41906 28700 41916 28756
rect 41972 28700 43484 28756
rect 43540 28700 43550 28756
rect 46498 28700 46508 28756
rect 46564 28700 47068 28756
rect 47124 28700 47162 28756
rect 29596 28644 29652 28700
rect 2594 28588 2604 28644
rect 2660 28588 3276 28644
rect 3332 28588 11340 28644
rect 11396 28588 11900 28644
rect 11956 28588 15148 28644
rect 17266 28588 17276 28644
rect 17332 28588 17836 28644
rect 17892 28588 17902 28644
rect 24882 28588 24892 28644
rect 24948 28588 25340 28644
rect 25396 28588 25564 28644
rect 25620 28588 25630 28644
rect 26450 28588 26460 28644
rect 26516 28588 29652 28644
rect 36642 28588 36652 28644
rect 36708 28588 42924 28644
rect 42980 28588 42990 28644
rect 44594 28588 44604 28644
rect 44660 28588 45052 28644
rect 45108 28588 48076 28644
rect 48132 28588 50428 28644
rect 50484 28588 50494 28644
rect 23426 28476 23436 28532
rect 23492 28476 23996 28532
rect 24052 28476 24062 28532
rect 28690 28476 28700 28532
rect 28756 28476 29036 28532
rect 29092 28476 29102 28532
rect 30258 28476 30268 28532
rect 30324 28476 30604 28532
rect 30660 28476 31052 28532
rect 31108 28476 34188 28532
rect 34244 28476 34254 28532
rect 36418 28476 36428 28532
rect 36484 28476 43372 28532
rect 43428 28476 43438 28532
rect 47170 28476 47180 28532
rect 47236 28476 47740 28532
rect 47796 28476 47806 28532
rect 6178 28364 6188 28420
rect 6244 28364 8988 28420
rect 9044 28364 9054 28420
rect 21970 28364 21980 28420
rect 22036 28364 25676 28420
rect 25732 28364 25742 28420
rect 29474 28364 29484 28420
rect 29540 28364 30044 28420
rect 30100 28364 30110 28420
rect 30370 28364 30380 28420
rect 30436 28364 30940 28420
rect 30996 28364 34076 28420
rect 34132 28364 34142 28420
rect 34738 28364 34748 28420
rect 34804 28364 43260 28420
rect 43316 28364 43326 28420
rect 40226 28252 40236 28308
rect 40292 28252 49532 28308
rect 49588 28252 49598 28308
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 50546 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50830 28252
rect 11554 28028 11564 28084
rect 11620 28028 12684 28084
rect 12740 28028 12750 28084
rect 16594 28028 16604 28084
rect 16660 28028 18844 28084
rect 18900 28028 18910 28084
rect 20514 28028 20524 28084
rect 20580 28028 22204 28084
rect 22260 28028 22270 28084
rect 23986 28028 23996 28084
rect 24052 28028 28252 28084
rect 28308 28028 28318 28084
rect 36418 28028 36428 28084
rect 36484 28028 37436 28084
rect 37492 28028 37502 28084
rect 41346 28028 41356 28084
rect 41412 28028 41804 28084
rect 41860 28028 41870 28084
rect 47394 28028 47404 28084
rect 47460 28028 48300 28084
rect 48356 28028 48972 28084
rect 49028 28028 49038 28084
rect 5618 27916 5628 27972
rect 5684 27916 5694 27972
rect 8194 27916 8204 27972
rect 8260 27916 11004 27972
rect 11060 27916 11070 27972
rect 15474 27916 15484 27972
rect 15540 27916 17500 27972
rect 17556 27916 17566 27972
rect 18386 27916 18396 27972
rect 18452 27916 19964 27972
rect 20020 27916 20030 27972
rect 21970 27916 21980 27972
rect 22036 27916 23772 27972
rect 23828 27916 23838 27972
rect 25442 27916 25452 27972
rect 25508 27916 31836 27972
rect 31892 27916 34860 27972
rect 34916 27916 37884 27972
rect 37940 27916 37950 27972
rect 5628 27860 5684 27916
rect 4946 27804 4956 27860
rect 5012 27804 6412 27860
rect 6468 27804 7420 27860
rect 7476 27804 16156 27860
rect 16212 27804 16222 27860
rect 16706 27804 16716 27860
rect 16772 27804 17164 27860
rect 17220 27804 17230 27860
rect 23426 27804 23436 27860
rect 23492 27748 23548 27860
rect 34738 27804 34748 27860
rect 34804 27804 35196 27860
rect 35252 27804 36092 27860
rect 36148 27804 36158 27860
rect 36754 27804 36764 27860
rect 36820 27804 37660 27860
rect 37716 27804 37726 27860
rect 16818 27692 16828 27748
rect 16884 27692 19404 27748
rect 19460 27692 19470 27748
rect 19618 27692 19628 27748
rect 19684 27692 19722 27748
rect 23492 27692 24220 27748
rect 24276 27692 24286 27748
rect 36306 27692 36316 27748
rect 36372 27692 37212 27748
rect 37268 27692 37278 27748
rect 43698 27692 43708 27748
rect 43764 27692 45276 27748
rect 45332 27692 45500 27748
rect 45556 27692 45566 27748
rect 17154 27580 17164 27636
rect 17220 27580 22428 27636
rect 22484 27580 22494 27636
rect 27458 27580 27468 27636
rect 27524 27580 39788 27636
rect 39844 27580 39854 27636
rect 19478 27468 19516 27524
rect 19572 27468 22204 27524
rect 22260 27468 22540 27524
rect 22596 27468 22606 27524
rect 28578 27468 28588 27524
rect 28644 27468 34748 27524
rect 34804 27468 34814 27524
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 54200 27412 55000 27440
rect 19282 27356 19292 27412
rect 19348 27356 28700 27412
rect 28756 27356 29708 27412
rect 29764 27356 29774 27412
rect 52658 27356 52668 27412
rect 52724 27356 53228 27412
rect 53284 27356 55000 27412
rect 54200 27328 55000 27356
rect 6178 27244 6188 27300
rect 6244 27244 6748 27300
rect 6804 27244 6814 27300
rect 24658 27244 24668 27300
rect 24724 27244 41356 27300
rect 41412 27244 41422 27300
rect 11554 27132 11564 27188
rect 11620 27132 11788 27188
rect 11844 27132 27468 27188
rect 27524 27132 27534 27188
rect 30594 27132 30604 27188
rect 30660 27132 31836 27188
rect 31892 27132 31902 27188
rect 35298 27132 35308 27188
rect 35364 27132 36652 27188
rect 36708 27132 36718 27188
rect 39778 27132 39788 27188
rect 39844 27132 45500 27188
rect 45556 27132 45566 27188
rect 8978 27020 8988 27076
rect 9044 27020 9772 27076
rect 9828 27020 11116 27076
rect 11172 27020 14700 27076
rect 14756 27020 14766 27076
rect 19058 27020 19068 27076
rect 19124 27020 19964 27076
rect 20020 27020 20030 27076
rect 22194 27020 22204 27076
rect 22260 27020 25004 27076
rect 25060 27020 25070 27076
rect 25666 27020 25676 27076
rect 25732 27020 26908 27076
rect 26852 26964 26908 27020
rect 29484 27020 30940 27076
rect 30996 27020 31006 27076
rect 33730 27020 33740 27076
rect 33796 27020 35756 27076
rect 35812 27020 35822 27076
rect 37762 27020 37772 27076
rect 37828 27020 41468 27076
rect 41524 27020 41534 27076
rect 43026 27020 43036 27076
rect 43092 27020 44156 27076
rect 44212 27020 44222 27076
rect 8866 26908 8876 26964
rect 8932 26908 9996 26964
rect 10052 26908 10780 26964
rect 10836 26908 10846 26964
rect 11666 26908 11676 26964
rect 11732 26908 12236 26964
rect 12292 26908 12302 26964
rect 19394 26908 19404 26964
rect 19460 26908 20300 26964
rect 20356 26908 20366 26964
rect 25218 26908 25228 26964
rect 25284 26908 26460 26964
rect 26516 26908 26526 26964
rect 26852 26908 28588 26964
rect 28644 26908 29260 26964
rect 29316 26908 29326 26964
rect 29484 26852 29540 27020
rect 30258 26908 30268 26964
rect 30324 26908 34076 26964
rect 34132 26908 34142 26964
rect 36082 26908 36092 26964
rect 36148 26908 39900 26964
rect 39956 26908 39966 26964
rect 42018 26908 42028 26964
rect 42084 26908 43708 26964
rect 43764 26908 43774 26964
rect 49634 26908 49644 26964
rect 49700 26908 50876 26964
rect 50932 26908 50942 26964
rect 23538 26796 23548 26852
rect 23604 26796 24108 26852
rect 24164 26796 24174 26852
rect 25330 26796 25340 26852
rect 25396 26796 25788 26852
rect 25844 26796 25854 26852
rect 29362 26796 29372 26852
rect 29428 26796 29540 26852
rect 29922 26796 29932 26852
rect 29988 26796 31724 26852
rect 31780 26796 31790 26852
rect 36530 26796 36540 26852
rect 36596 26796 37996 26852
rect 38052 26796 38062 26852
rect 29698 26684 29708 26740
rect 29764 26684 30268 26740
rect 30324 26684 30334 26740
rect 31490 26684 31500 26740
rect 31556 26684 33964 26740
rect 34020 26684 35308 26740
rect 35364 26684 35980 26740
rect 36036 26684 36046 26740
rect 39442 26684 39452 26740
rect 39508 26684 40124 26740
rect 40180 26684 40190 26740
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 50546 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50830 26684
rect 28802 26572 28812 26628
rect 28868 26572 29260 26628
rect 29316 26572 31164 26628
rect 31220 26572 33852 26628
rect 33908 26572 34748 26628
rect 34804 26572 34814 26628
rect 35186 26572 35196 26628
rect 35252 26572 35756 26628
rect 35812 26572 35822 26628
rect 2482 26460 2492 26516
rect 2548 26460 3388 26516
rect 5954 26460 5964 26516
rect 6020 26460 7756 26516
rect 7812 26460 7822 26516
rect 26226 26460 26236 26516
rect 26292 26460 42364 26516
rect 42420 26460 42430 26516
rect 3332 26180 3388 26460
rect 28914 26348 28924 26404
rect 28980 26348 30828 26404
rect 30884 26348 31500 26404
rect 31556 26348 31566 26404
rect 8418 26236 8428 26292
rect 8484 26236 9548 26292
rect 9604 26236 9614 26292
rect 33506 26236 33516 26292
rect 33572 26236 38780 26292
rect 38836 26236 38846 26292
rect 3332 26124 5404 26180
rect 5460 26124 5470 26180
rect 28018 26124 28028 26180
rect 28084 26124 29484 26180
rect 29540 26124 29550 26180
rect 30258 26124 30268 26180
rect 30324 26124 37324 26180
rect 37380 26124 37390 26180
rect 41346 26124 41356 26180
rect 41412 26124 42140 26180
rect 42196 26124 42924 26180
rect 42980 26124 42990 26180
rect 49522 26124 49532 26180
rect 49588 26124 50988 26180
rect 51044 26124 51054 26180
rect 38882 26012 38892 26068
rect 38948 26012 39676 26068
rect 39732 26012 39742 26068
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 37986 25788 37996 25844
rect 38052 25788 39340 25844
rect 39396 25788 39406 25844
rect 7746 25676 7756 25732
rect 7812 25676 7822 25732
rect 7970 25676 7980 25732
rect 8036 25676 8540 25732
rect 8596 25676 8606 25732
rect 31892 25676 38668 25732
rect 38724 25676 38734 25732
rect 7756 25620 7812 25676
rect 31892 25620 31948 25676
rect 7756 25564 8932 25620
rect 15138 25564 15148 25620
rect 15204 25564 17724 25620
rect 17780 25564 17790 25620
rect 26338 25564 26348 25620
rect 26404 25564 31948 25620
rect 32050 25564 32060 25620
rect 32116 25564 33628 25620
rect 33684 25564 33694 25620
rect 36194 25564 36204 25620
rect 36260 25564 37156 25620
rect 37314 25564 37324 25620
rect 37380 25564 38668 25620
rect 50082 25564 50092 25620
rect 50148 25564 53228 25620
rect 53284 25564 53294 25620
rect 8876 25396 8932 25564
rect 37100 25508 37156 25564
rect 38612 25508 38668 25564
rect 9650 25452 9660 25508
rect 9716 25452 11116 25508
rect 11172 25452 11182 25508
rect 19506 25452 19516 25508
rect 19572 25452 19852 25508
rect 19908 25452 19918 25508
rect 23874 25452 23884 25508
rect 23940 25452 24556 25508
rect 24612 25452 25788 25508
rect 25844 25452 25854 25508
rect 30034 25452 30044 25508
rect 30100 25452 35420 25508
rect 35476 25452 36316 25508
rect 36372 25452 36382 25508
rect 37090 25452 37100 25508
rect 37156 25452 38108 25508
rect 38164 25452 38174 25508
rect 38612 25452 40852 25508
rect 46050 25452 46060 25508
rect 46116 25452 47740 25508
rect 47796 25452 49420 25508
rect 49476 25452 49486 25508
rect 40796 25396 40852 25452
rect 4386 25340 4396 25396
rect 4452 25340 7196 25396
rect 7252 25340 8204 25396
rect 8260 25340 8652 25396
rect 8708 25340 8718 25396
rect 8876 25340 9828 25396
rect 16818 25340 16828 25396
rect 16884 25340 17612 25396
rect 17668 25340 17678 25396
rect 24098 25340 24108 25396
rect 24164 25340 25228 25396
rect 25284 25340 25294 25396
rect 29810 25340 29820 25396
rect 29876 25340 31164 25396
rect 31220 25340 31836 25396
rect 31892 25340 32228 25396
rect 39330 25340 39340 25396
rect 39396 25340 39900 25396
rect 39956 25340 39966 25396
rect 40786 25340 40796 25396
rect 40852 25340 40862 25396
rect 46162 25340 46172 25396
rect 46228 25340 47964 25396
rect 48020 25340 48188 25396
rect 48244 25340 48254 25396
rect 49298 25340 49308 25396
rect 49364 25340 50204 25396
rect 50260 25340 50270 25396
rect 6402 25228 6412 25284
rect 6468 25228 7308 25284
rect 7364 25228 8428 25284
rect 8484 25228 8494 25284
rect 9772 25060 9828 25340
rect 32172 25284 32228 25340
rect 10994 25228 11004 25284
rect 11060 25228 11900 25284
rect 11956 25228 11966 25284
rect 17714 25228 17724 25284
rect 17780 25228 19740 25284
rect 19796 25228 20300 25284
rect 20356 25228 22988 25284
rect 23044 25228 23054 25284
rect 29708 25228 30380 25284
rect 30436 25228 31892 25284
rect 31948 25228 31958 25284
rect 32172 25228 37324 25284
rect 37380 25228 37390 25284
rect 37538 25228 37548 25284
rect 37604 25228 38556 25284
rect 38612 25228 42252 25284
rect 42308 25228 42318 25284
rect 48402 25228 48412 25284
rect 48468 25228 48860 25284
rect 48916 25228 48926 25284
rect 29708 25172 29764 25228
rect 37548 25172 37604 25228
rect 20514 25116 20524 25172
rect 20580 25116 21084 25172
rect 21140 25116 29708 25172
rect 29764 25116 29774 25172
rect 32274 25116 32284 25172
rect 32340 25116 37604 25172
rect 40226 25116 40236 25172
rect 40292 25116 46396 25172
rect 46452 25116 46462 25172
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 50546 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50830 25116
rect 9762 25004 9772 25060
rect 9828 25004 9838 25060
rect 29026 25004 29036 25060
rect 29092 25004 37660 25060
rect 37716 25004 37726 25060
rect 43138 25004 43148 25060
rect 43204 25004 44044 25060
rect 44100 25004 44110 25060
rect 11106 24892 11116 24948
rect 11172 24892 11900 24948
rect 11956 24892 11966 24948
rect 16706 24892 16716 24948
rect 16772 24892 17500 24948
rect 17556 24892 21868 24948
rect 21924 24892 22316 24948
rect 22372 24892 24668 24948
rect 24724 24892 25564 24948
rect 25620 24892 25630 24948
rect 25778 24892 25788 24948
rect 25844 24892 26796 24948
rect 26852 24892 26862 24948
rect 29138 24892 29148 24948
rect 29204 24892 33516 24948
rect 33572 24892 33582 24948
rect 39442 24892 39452 24948
rect 39508 24892 39788 24948
rect 39844 24892 39854 24948
rect 4722 24780 4732 24836
rect 4788 24780 5404 24836
rect 5460 24780 7644 24836
rect 7700 24780 7710 24836
rect 20626 24780 20636 24836
rect 20692 24780 22988 24836
rect 23044 24780 23054 24836
rect 31378 24780 31388 24836
rect 31444 24780 32284 24836
rect 32340 24780 32350 24836
rect 54200 24724 55000 24752
rect 10658 24668 10668 24724
rect 10724 24668 11564 24724
rect 11620 24668 14476 24724
rect 14532 24668 16156 24724
rect 16212 24668 16222 24724
rect 19842 24668 19852 24724
rect 19908 24668 20300 24724
rect 20356 24668 20366 24724
rect 26226 24668 26236 24724
rect 26292 24668 28812 24724
rect 28868 24668 28878 24724
rect 31154 24668 31164 24724
rect 31220 24668 32172 24724
rect 32228 24668 32238 24724
rect 33842 24668 33852 24724
rect 33908 24668 37100 24724
rect 37156 24668 37166 24724
rect 37762 24668 37772 24724
rect 37828 24668 38556 24724
rect 38612 24668 41076 24724
rect 42242 24668 42252 24724
rect 42308 24668 43484 24724
rect 43540 24668 43550 24724
rect 53218 24668 53228 24724
rect 53284 24668 55000 24724
rect 5170 24556 5180 24612
rect 5236 24556 10108 24612
rect 10164 24556 11116 24612
rect 11172 24556 11676 24612
rect 11732 24556 12348 24612
rect 12404 24556 12414 24612
rect 39638 24556 39676 24612
rect 39732 24556 39742 24612
rect 41020 24500 41076 24668
rect 54200 24640 55000 24668
rect 41234 24556 41244 24612
rect 41300 24556 43148 24612
rect 43204 24556 43214 24612
rect 49074 24556 49084 24612
rect 49140 24556 49644 24612
rect 49700 24556 50204 24612
rect 50260 24556 50652 24612
rect 50708 24556 50718 24612
rect 31266 24444 31276 24500
rect 31332 24444 32172 24500
rect 32228 24444 32238 24500
rect 33282 24444 33292 24500
rect 33348 24444 34188 24500
rect 34244 24444 34254 24500
rect 34850 24444 34860 24500
rect 34916 24444 36652 24500
rect 36708 24444 40012 24500
rect 40068 24444 40078 24500
rect 41020 24444 42140 24500
rect 42196 24444 42206 24500
rect 18386 24332 18396 24388
rect 18452 24332 19292 24388
rect 19348 24332 29932 24388
rect 29988 24332 29998 24388
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 6066 24220 6076 24276
rect 6132 24220 6142 24276
rect 6076 24164 6132 24220
rect 4498 24108 4508 24164
rect 4564 24108 6132 24164
rect 35186 24108 35196 24164
rect 35252 24108 36988 24164
rect 37044 24108 37054 24164
rect 26114 23996 26124 24052
rect 26180 23996 33404 24052
rect 33460 23996 33470 24052
rect 36204 23996 47068 24052
rect 47124 23996 47134 24052
rect 49420 23996 52556 24052
rect 52612 23996 52622 24052
rect 8194 23884 8204 23940
rect 8260 23884 8540 23940
rect 8596 23884 8876 23940
rect 8932 23884 15148 23940
rect 15698 23884 15708 23940
rect 15764 23884 18060 23940
rect 18116 23884 18126 23940
rect 15092 23828 15148 23884
rect 6066 23772 6076 23828
rect 6132 23772 8764 23828
rect 8820 23772 10556 23828
rect 10612 23772 10622 23828
rect 15092 23772 15372 23828
rect 15428 23772 15438 23828
rect 2818 23660 2828 23716
rect 2884 23660 5964 23716
rect 6020 23660 6030 23716
rect 8306 23660 8316 23716
rect 8372 23660 9100 23716
rect 9156 23660 9166 23716
rect 20066 23660 20076 23716
rect 20132 23660 21420 23716
rect 21476 23660 21486 23716
rect 25218 23660 25228 23716
rect 25284 23660 26124 23716
rect 26180 23660 26190 23716
rect 30930 23660 30940 23716
rect 30996 23660 34972 23716
rect 35028 23660 35038 23716
rect 36204 23604 36260 23996
rect 37650 23884 37660 23940
rect 37716 23884 39564 23940
rect 39620 23884 39630 23940
rect 46162 23884 46172 23940
rect 46228 23884 46238 23940
rect 37986 23772 37996 23828
rect 38052 23772 38780 23828
rect 38836 23772 38846 23828
rect 43586 23772 43596 23828
rect 43652 23772 44044 23828
rect 44100 23772 44828 23828
rect 44884 23772 44894 23828
rect 46172 23716 46228 23884
rect 49420 23716 49476 23996
rect 49644 23884 52892 23940
rect 52948 23884 52958 23940
rect 37314 23660 37324 23716
rect 37380 23660 46228 23716
rect 47618 23660 47628 23716
rect 47684 23660 49420 23716
rect 49476 23660 49486 23716
rect 49644 23604 49700 23884
rect 1810 23548 1820 23604
rect 1876 23548 5068 23604
rect 5124 23548 5516 23604
rect 5572 23548 5582 23604
rect 33618 23548 33628 23604
rect 33684 23548 34636 23604
rect 34692 23548 36260 23604
rect 40348 23548 44604 23604
rect 44660 23548 44670 23604
rect 45714 23548 45724 23604
rect 45780 23548 45790 23604
rect 46722 23548 46732 23604
rect 46788 23548 48300 23604
rect 48356 23548 49700 23604
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 40348 23492 40404 23548
rect 45724 23492 45780 23548
rect 50546 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50830 23548
rect 4946 23436 4956 23492
rect 5012 23436 5852 23492
rect 5908 23436 6524 23492
rect 6580 23436 7196 23492
rect 7252 23436 7262 23492
rect 20626 23436 20636 23492
rect 20692 23436 22092 23492
rect 22148 23436 22158 23492
rect 25666 23436 25676 23492
rect 25732 23436 26684 23492
rect 26740 23436 26750 23492
rect 39442 23436 39452 23492
rect 39508 23436 40404 23492
rect 42578 23436 42588 23492
rect 42644 23436 43596 23492
rect 43652 23436 43662 23492
rect 45378 23436 45388 23492
rect 45444 23436 46620 23492
rect 46676 23436 46686 23492
rect 5394 23324 5404 23380
rect 5460 23324 6468 23380
rect 28018 23324 28028 23380
rect 28084 23324 31500 23380
rect 31556 23324 31566 23380
rect 43250 23324 43260 23380
rect 43316 23324 43326 23380
rect 45602 23324 45612 23380
rect 45668 23324 46172 23380
rect 46228 23324 46396 23380
rect 46452 23324 46462 23380
rect 6412 23268 6468 23324
rect 4946 23212 4956 23268
rect 5012 23212 6188 23268
rect 6244 23212 6254 23268
rect 6402 23212 6412 23268
rect 6468 23212 7644 23268
rect 7700 23212 7710 23268
rect 36642 23100 36652 23156
rect 36708 23100 40012 23156
rect 40068 23100 40078 23156
rect 43260 23044 43316 23324
rect 50372 23156 50428 23268
rect 50484 23212 50494 23268
rect 43474 23100 43484 23156
rect 43540 23100 44156 23156
rect 44212 23100 44222 23156
rect 47964 23100 50428 23156
rect 47964 23044 48020 23100
rect 7410 22988 7420 23044
rect 7476 22988 8428 23044
rect 8484 22988 8494 23044
rect 8978 22988 8988 23044
rect 9044 22988 13468 23044
rect 13524 22988 13534 23044
rect 29362 22988 29372 23044
rect 29428 22988 30380 23044
rect 30436 22988 36428 23044
rect 36484 22988 36494 23044
rect 37202 22988 37212 23044
rect 37268 22988 37548 23044
rect 37604 22988 38444 23044
rect 38500 22988 38510 23044
rect 42130 22988 42140 23044
rect 42196 22988 42700 23044
rect 42756 22988 42766 23044
rect 42914 22988 42924 23044
rect 42980 22988 44492 23044
rect 44548 22988 44558 23044
rect 47954 22988 47964 23044
rect 48020 22988 48030 23044
rect 49522 22988 49532 23044
rect 49588 22988 50876 23044
rect 50932 22988 50942 23044
rect 5058 22876 5068 22932
rect 5124 22876 5628 22932
rect 5684 22876 5694 22932
rect 8866 22876 8876 22932
rect 8932 22876 9212 22932
rect 9268 22876 20636 22932
rect 20692 22876 20702 22932
rect 26898 22876 26908 22932
rect 26964 22876 42588 22932
rect 42644 22876 42654 22932
rect 46274 22876 46284 22932
rect 46340 22876 49308 22932
rect 49364 22876 49374 22932
rect 41346 22764 41356 22820
rect 41412 22764 43260 22820
rect 43316 22764 43326 22820
rect 50082 22764 50092 22820
rect 50148 22764 50316 22820
rect 50372 22764 50382 22820
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 26674 22428 26684 22484
rect 26740 22428 48916 22484
rect 50418 22428 50428 22484
rect 50484 22428 53228 22484
rect 53284 22428 53294 22484
rect 21746 22316 21756 22372
rect 21812 22316 21822 22372
rect 23650 22316 23660 22372
rect 23716 22316 24332 22372
rect 24388 22316 24398 22372
rect 5926 22204 5964 22260
rect 6020 22204 6636 22260
rect 6692 22204 6702 22260
rect 21756 22148 21812 22316
rect 26852 22260 26908 22428
rect 28242 22316 28252 22372
rect 28308 22316 29148 22372
rect 29204 22316 29214 22372
rect 33954 22316 33964 22372
rect 34020 22316 36988 22372
rect 37044 22316 37054 22372
rect 39218 22316 39228 22372
rect 39284 22316 40012 22372
rect 40068 22316 41244 22372
rect 41300 22316 41310 22372
rect 42690 22316 42700 22372
rect 42756 22316 43484 22372
rect 43540 22316 43550 22372
rect 26450 22204 26460 22260
rect 26516 22204 26908 22260
rect 29474 22204 29484 22260
rect 29540 22204 30828 22260
rect 30884 22204 30894 22260
rect 35410 22204 35420 22260
rect 35476 22204 37324 22260
rect 37380 22204 37390 22260
rect 37772 22204 38668 22260
rect 41430 22204 41468 22260
rect 41524 22204 41534 22260
rect 45378 22204 45388 22260
rect 45444 22204 46284 22260
rect 46340 22204 46350 22260
rect 2482 22092 2492 22148
rect 2548 22092 5740 22148
rect 5796 22092 5806 22148
rect 20402 22092 20412 22148
rect 20468 22092 23996 22148
rect 24052 22092 24062 22148
rect 25890 22092 25900 22148
rect 25956 22092 25966 22148
rect 26562 22092 26572 22148
rect 26628 22092 34860 22148
rect 34916 22092 35308 22148
rect 35364 22092 35374 22148
rect 25900 22036 25956 22092
rect 37772 22036 37828 22204
rect 25900 21980 26908 22036
rect 26964 21980 37828 22036
rect 38612 22036 38668 22204
rect 48860 22148 48916 22428
rect 49746 22204 49756 22260
rect 49812 22204 50204 22260
rect 50260 22204 50270 22260
rect 40450 22092 40460 22148
rect 40516 22092 41692 22148
rect 41748 22092 42364 22148
rect 42420 22092 42430 22148
rect 42690 22092 42700 22148
rect 42756 22092 43820 22148
rect 43876 22092 44268 22148
rect 44324 22092 44492 22148
rect 44548 22092 44558 22148
rect 45042 22092 45052 22148
rect 45108 22092 47852 22148
rect 47908 22092 47918 22148
rect 48850 22092 48860 22148
rect 48916 22092 50036 22148
rect 49980 22036 50036 22092
rect 54200 22036 55000 22064
rect 38612 21980 46620 22036
rect 46676 21980 46686 22036
rect 49942 21980 49980 22036
rect 50036 21980 50046 22036
rect 53330 21980 53340 22036
rect 53396 21980 55000 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 50546 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50830 21980
rect 54200 21952 55000 21980
rect 9986 21868 9996 21924
rect 10052 21868 10062 21924
rect 24658 21868 24668 21924
rect 24724 21868 25564 21924
rect 25620 21868 26348 21924
rect 26404 21868 26414 21924
rect 30818 21868 30828 21924
rect 30884 21868 33964 21924
rect 34020 21868 34030 21924
rect 37538 21868 37548 21924
rect 37604 21868 40908 21924
rect 40964 21868 41356 21924
rect 41412 21868 41422 21924
rect 41580 21868 45388 21924
rect 45444 21868 45454 21924
rect 49858 21868 49868 21924
rect 49924 21868 50092 21924
rect 50148 21868 50158 21924
rect 9996 21812 10052 21868
rect 4610 21756 4620 21812
rect 4676 21756 5292 21812
rect 5348 21756 5358 21812
rect 8082 21756 8092 21812
rect 8148 21756 8652 21812
rect 8708 21756 8718 21812
rect 9650 21756 9660 21812
rect 9716 21756 10052 21812
rect 12674 21756 12684 21812
rect 12740 21756 14028 21812
rect 14084 21756 14094 21812
rect 21858 21756 21868 21812
rect 21924 21756 22204 21812
rect 22260 21756 22652 21812
rect 22708 21756 23548 21812
rect 23604 21756 23614 21812
rect 35298 21756 35308 21812
rect 35364 21756 37212 21812
rect 37268 21756 38556 21812
rect 38612 21756 38622 21812
rect 9996 21700 10052 21756
rect 41580 21700 41636 21868
rect 42802 21756 42812 21812
rect 42868 21756 43596 21812
rect 43652 21756 43662 21812
rect 46386 21756 46396 21812
rect 46452 21756 49420 21812
rect 49476 21756 52892 21812
rect 52948 21756 52958 21812
rect 9996 21644 11340 21700
rect 11396 21644 13468 21700
rect 13524 21644 16940 21700
rect 16996 21644 17006 21700
rect 22978 21644 22988 21700
rect 23044 21644 23884 21700
rect 23940 21644 27020 21700
rect 27076 21644 27692 21700
rect 27748 21644 27758 21700
rect 30594 21644 30604 21700
rect 30660 21644 30940 21700
rect 30996 21644 33180 21700
rect 33236 21644 33246 21700
rect 37986 21644 37996 21700
rect 38052 21644 39228 21700
rect 39284 21644 40348 21700
rect 40404 21644 41580 21700
rect 41636 21644 41646 21700
rect 43026 21644 43036 21700
rect 43092 21644 43484 21700
rect 43540 21644 43550 21700
rect 47954 21644 47964 21700
rect 48020 21644 48748 21700
rect 48804 21644 49308 21700
rect 49364 21644 49374 21700
rect 9996 21476 10052 21644
rect 23202 21532 23212 21588
rect 23268 21532 24780 21588
rect 24836 21532 24846 21588
rect 30818 21532 30828 21588
rect 30884 21532 31612 21588
rect 31668 21532 38668 21588
rect 40226 21532 40236 21588
rect 40292 21532 41132 21588
rect 41188 21532 41198 21588
rect 43922 21532 43932 21588
rect 43988 21532 45276 21588
rect 45332 21532 45342 21588
rect 45826 21532 45836 21588
rect 45892 21532 45902 21588
rect 47282 21532 47292 21588
rect 47348 21532 48636 21588
rect 48692 21532 52780 21588
rect 52836 21532 52846 21588
rect 38612 21476 38668 21532
rect 45836 21476 45892 21532
rect 9986 21420 9996 21476
rect 10052 21420 10062 21476
rect 31714 21420 31724 21476
rect 31780 21420 33404 21476
rect 33460 21420 33470 21476
rect 37090 21420 37100 21476
rect 37156 21420 37660 21476
rect 37716 21420 38108 21476
rect 38164 21420 38174 21476
rect 38612 21420 45892 21476
rect 15026 21308 15036 21364
rect 15092 21308 21532 21364
rect 21588 21308 22316 21364
rect 22372 21308 31948 21364
rect 41234 21308 41244 21364
rect 41300 21308 42812 21364
rect 42868 21308 42878 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 31892 21028 31948 21308
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 38612 21084 41020 21140
rect 41076 21084 41086 21140
rect 38612 21028 38668 21084
rect 9874 20972 9884 21028
rect 9940 20972 10556 21028
rect 10612 20972 10622 21028
rect 31892 20972 38668 21028
rect 45714 20972 45724 21028
rect 45780 20972 46508 21028
rect 46564 20972 46574 21028
rect 18498 20860 18508 20916
rect 18564 20860 37548 20916
rect 37604 20860 37614 20916
rect 48066 20860 48076 20916
rect 48132 20860 49980 20916
rect 50036 20860 50046 20916
rect 10966 20748 11004 20804
rect 11060 20748 11070 20804
rect 27010 20748 27020 20804
rect 27076 20748 27916 20804
rect 27972 20748 27982 20804
rect 28466 20748 28476 20804
rect 28532 20748 30268 20804
rect 30324 20748 30334 20804
rect 32050 20748 32060 20804
rect 32116 20748 45948 20804
rect 46004 20748 46014 20804
rect 46498 20748 46508 20804
rect 46564 20748 48860 20804
rect 48916 20748 52892 20804
rect 52948 20748 52958 20804
rect 8754 20636 8764 20692
rect 8820 20636 13804 20692
rect 13860 20636 15260 20692
rect 15316 20636 16380 20692
rect 16436 20636 16446 20692
rect 16706 20636 16716 20692
rect 16772 20636 18844 20692
rect 18900 20636 18910 20692
rect 19058 20636 19068 20692
rect 19124 20636 19628 20692
rect 19684 20636 19694 20692
rect 27682 20636 27692 20692
rect 27748 20636 29036 20692
rect 29092 20636 29102 20692
rect 44930 20636 44940 20692
rect 44996 20636 45892 20692
rect 45836 20580 45892 20636
rect 18284 20524 39564 20580
rect 39620 20524 39630 20580
rect 45826 20524 45836 20580
rect 45892 20524 46956 20580
rect 47012 20524 47022 20580
rect 18284 20468 18340 20524
rect 8642 20412 8652 20468
rect 8708 20412 9660 20468
rect 9716 20412 18340 20468
rect 27906 20412 27916 20468
rect 27972 20412 28364 20468
rect 28420 20412 28430 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 50546 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50830 20412
rect 20962 20188 20972 20244
rect 21028 20188 22204 20244
rect 22260 20188 22270 20244
rect 30034 20188 30044 20244
rect 30100 20188 30492 20244
rect 30548 20188 30558 20244
rect 39554 20188 39564 20244
rect 39620 20188 40124 20244
rect 40180 20188 40190 20244
rect 43222 20188 43260 20244
rect 43316 20188 44156 20244
rect 44212 20188 44222 20244
rect 45490 20188 45500 20244
rect 45556 20188 46396 20244
rect 46452 20188 47404 20244
rect 47460 20188 47628 20244
rect 47684 20188 47694 20244
rect 7074 20076 7084 20132
rect 7140 20076 8652 20132
rect 8708 20076 8718 20132
rect 14466 20076 14476 20132
rect 14532 20076 15820 20132
rect 15876 20076 15886 20132
rect 16482 20076 16492 20132
rect 16548 20076 16558 20132
rect 24770 20076 24780 20132
rect 24836 20076 25788 20132
rect 25844 20076 25854 20132
rect 27234 20076 27244 20132
rect 27300 20076 28476 20132
rect 28532 20076 28542 20132
rect 8306 19964 8316 20020
rect 8372 19964 8988 20020
rect 9044 19964 9054 20020
rect 14914 19964 14924 20020
rect 14980 19964 15484 20020
rect 15540 19964 16156 20020
rect 16212 19964 16222 20020
rect 16492 19908 16548 20076
rect 25526 19964 25564 20020
rect 25620 19964 25630 20020
rect 28018 19964 28028 20020
rect 28084 19964 28812 20020
rect 28868 19964 28878 20020
rect 4946 19852 4956 19908
rect 5012 19852 6412 19908
rect 6468 19852 9772 19908
rect 9828 19852 9838 19908
rect 12002 19852 12012 19908
rect 12068 19852 16548 19908
rect 23986 19852 23996 19908
rect 24052 19852 25340 19908
rect 25396 19852 25406 19908
rect 28130 19852 28140 19908
rect 28196 19852 31612 19908
rect 31668 19852 31678 19908
rect 40898 19852 40908 19908
rect 40964 19852 45948 19908
rect 46004 19852 46014 19908
rect 50194 19852 50204 19908
rect 50260 19852 53228 19908
rect 53284 19852 53294 19908
rect 7074 19740 7084 19796
rect 7140 19740 7644 19796
rect 7700 19740 8876 19796
rect 8932 19740 8942 19796
rect 10098 19740 10108 19796
rect 10164 19740 11116 19796
rect 11172 19740 15148 19796
rect 15204 19740 15214 19796
rect 16594 19740 16604 19796
rect 16660 19740 39788 19796
rect 39844 19740 39854 19796
rect 46050 19740 46060 19796
rect 46116 19740 46844 19796
rect 46900 19740 50540 19796
rect 50596 19740 50606 19796
rect 22082 19628 22092 19684
rect 22148 19628 23436 19684
rect 23492 19628 28700 19684
rect 28756 19628 29260 19684
rect 29316 19628 31052 19684
rect 31108 19628 31118 19684
rect 38966 19628 39004 19684
rect 39060 19628 39070 19684
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 39750 19516 39788 19572
rect 39844 19516 39854 19572
rect 8978 19404 8988 19460
rect 9044 19404 11452 19460
rect 11508 19404 17052 19460
rect 17108 19404 17118 19460
rect 31154 19404 31164 19460
rect 31220 19404 38444 19460
rect 38500 19404 38510 19460
rect 54200 19348 55000 19376
rect 7970 19292 7980 19348
rect 8036 19292 8540 19348
rect 8596 19292 9100 19348
rect 9156 19292 11228 19348
rect 11284 19292 12012 19348
rect 12068 19292 12078 19348
rect 32498 19292 32508 19348
rect 32564 19292 34300 19348
rect 34356 19292 34860 19348
rect 34916 19292 34926 19348
rect 53218 19292 53228 19348
rect 53284 19292 55000 19348
rect 54200 19264 55000 19292
rect 31164 19180 31612 19236
rect 31668 19180 32172 19236
rect 32228 19180 32238 19236
rect 33282 19180 33292 19236
rect 33348 19180 35308 19236
rect 35364 19180 35374 19236
rect 45602 19180 45612 19236
rect 45668 19180 45948 19236
rect 46004 19180 46284 19236
rect 46340 19180 46350 19236
rect 46610 19180 46620 19236
rect 46676 19180 50988 19236
rect 51044 19180 51054 19236
rect 31164 19124 31220 19180
rect 7074 19068 7084 19124
rect 7140 19068 8316 19124
rect 8372 19068 10108 19124
rect 10164 19068 14364 19124
rect 14420 19068 14430 19124
rect 31154 19068 31164 19124
rect 31220 19068 31230 19124
rect 31826 19068 31836 19124
rect 31892 19068 32844 19124
rect 32900 19068 32910 19124
rect 34626 19068 34636 19124
rect 34692 19068 35196 19124
rect 35252 19068 35262 19124
rect 47954 19068 47964 19124
rect 48020 19068 48412 19124
rect 48468 19068 48478 19124
rect 50194 19068 50204 19124
rect 50260 19068 50764 19124
rect 50820 19068 50830 19124
rect 4946 18956 4956 19012
rect 5012 18956 5628 19012
rect 5684 18956 5694 19012
rect 6178 18956 6188 19012
rect 6244 18956 10444 19012
rect 10500 18956 11004 19012
rect 11060 18956 11070 19012
rect 21522 18956 21532 19012
rect 21588 18956 22540 19012
rect 22596 18956 22606 19012
rect 30706 18956 30716 19012
rect 30772 18956 32620 19012
rect 32676 18956 32686 19012
rect 33954 18956 33964 19012
rect 34020 18956 34412 19012
rect 34468 18956 46732 19012
rect 46788 18956 46798 19012
rect 48178 18956 48188 19012
rect 48244 18956 50316 19012
rect 33964 18900 34020 18956
rect 6626 18844 6636 18900
rect 6692 18844 6702 18900
rect 30930 18844 30940 18900
rect 30996 18844 31276 18900
rect 31332 18844 34020 18900
rect 42130 18844 42140 18900
rect 42196 18844 43260 18900
rect 43316 18844 43372 18900
rect 43428 18844 43438 18900
rect 49298 18844 49308 18900
rect 49364 18844 50092 18900
rect 50148 18844 50158 18900
rect 6636 18452 6692 18844
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 50372 18676 50428 19012
rect 50546 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50830 18844
rect 38612 18620 39004 18676
rect 39060 18620 39070 18676
rect 50372 18620 50540 18676
rect 50596 18620 50606 18676
rect 38612 18564 38668 18620
rect 22866 18508 22876 18564
rect 22932 18508 23660 18564
rect 23716 18508 23726 18564
rect 25330 18508 25340 18564
rect 25396 18508 26012 18564
rect 26068 18508 26078 18564
rect 36418 18508 36428 18564
rect 36484 18508 38332 18564
rect 38388 18508 38668 18564
rect 39004 18564 39060 18620
rect 39004 18508 42028 18564
rect 42084 18508 42094 18564
rect 42578 18508 42588 18564
rect 42644 18508 45500 18564
rect 45556 18508 46172 18564
rect 46228 18508 46238 18564
rect 2482 18396 2492 18452
rect 2548 18396 6692 18452
rect 34962 18396 34972 18452
rect 35028 18396 36092 18452
rect 36148 18396 36158 18452
rect 38612 18396 38892 18452
rect 38948 18396 40348 18452
rect 40404 18396 41020 18452
rect 41076 18396 41804 18452
rect 41860 18396 42252 18452
rect 42308 18396 42318 18452
rect 45826 18396 45836 18452
rect 45892 18396 49196 18452
rect 49252 18396 49262 18452
rect 38612 18340 38668 18396
rect 4610 18284 4620 18340
rect 4676 18284 5516 18340
rect 5572 18284 5582 18340
rect 35410 18284 35420 18340
rect 35476 18284 38668 18340
rect 41906 18284 41916 18340
rect 41972 18284 42924 18340
rect 42980 18284 42990 18340
rect 43250 18284 43260 18340
rect 43316 18284 45052 18340
rect 45108 18284 45118 18340
rect 46162 18284 46172 18340
rect 46228 18284 46238 18340
rect 50306 18284 50316 18340
rect 50372 18284 50876 18340
rect 50932 18284 50942 18340
rect 46172 18228 46228 18284
rect 31042 18172 31052 18228
rect 31108 18172 46228 18228
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 48850 17836 48860 17892
rect 48916 17836 49756 17892
rect 49812 17836 49822 17892
rect 6402 17724 6412 17780
rect 6468 17724 6972 17780
rect 7028 17724 7980 17780
rect 8036 17724 8046 17780
rect 14802 17724 14812 17780
rect 14868 17724 15708 17780
rect 15764 17724 22092 17780
rect 22148 17724 22158 17780
rect 38546 17724 38556 17780
rect 38612 17724 39564 17780
rect 39620 17724 39630 17780
rect 21858 17612 21868 17668
rect 21924 17612 22876 17668
rect 22932 17612 22942 17668
rect 25890 17612 25900 17668
rect 25956 17612 29596 17668
rect 29652 17612 30044 17668
rect 30100 17612 30110 17668
rect 38098 17612 38108 17668
rect 38164 17612 40460 17668
rect 40516 17612 40526 17668
rect 48514 17612 48524 17668
rect 48580 17612 49308 17668
rect 49364 17612 49374 17668
rect 5506 17500 5516 17556
rect 5572 17500 6300 17556
rect 6356 17500 6366 17556
rect 14690 17500 14700 17556
rect 14756 17500 15148 17556
rect 15204 17500 15214 17556
rect 23650 17500 23660 17556
rect 23716 17500 25452 17556
rect 25508 17500 25518 17556
rect 32946 17500 32956 17556
rect 33012 17500 33404 17556
rect 33460 17500 34748 17556
rect 34804 17500 38556 17556
rect 38612 17500 38622 17556
rect 47618 17500 47628 17556
rect 47684 17500 48188 17556
rect 48244 17500 48254 17556
rect 32722 17388 32732 17444
rect 32788 17388 33516 17444
rect 33572 17388 33582 17444
rect 35074 17388 35084 17444
rect 35140 17388 36316 17444
rect 36372 17388 37884 17444
rect 37940 17388 37950 17444
rect 47170 17388 47180 17444
rect 47236 17388 47740 17444
rect 47796 17388 48860 17444
rect 48916 17388 52332 17444
rect 52388 17388 52398 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 50546 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50830 17276
rect 10546 17164 10556 17220
rect 10612 17164 13468 17220
rect 13524 17164 15148 17220
rect 11554 17052 11564 17108
rect 11620 17052 12348 17108
rect 12404 17052 12414 17108
rect 13122 17052 13132 17108
rect 13188 17052 14868 17108
rect 10210 16940 10220 16996
rect 10276 16940 11676 16996
rect 11732 16940 13020 16996
rect 13076 16940 13086 16996
rect 14812 16884 14868 17052
rect 15092 16996 15148 17164
rect 18162 17052 18172 17108
rect 18228 17052 19292 17108
rect 19348 17052 19358 17108
rect 32946 17052 32956 17108
rect 33012 17052 35308 17108
rect 35364 17052 35374 17108
rect 49186 17052 49196 17108
rect 49252 17052 49644 17108
rect 49700 17052 49710 17108
rect 15092 16940 16716 16996
rect 16772 16940 16782 16996
rect 32834 16940 32844 16996
rect 32900 16940 33404 16996
rect 33460 16940 33470 16996
rect 34178 16940 34188 16996
rect 34244 16940 35420 16996
rect 35476 16940 35486 16996
rect 42018 16940 42028 16996
rect 42084 16940 42700 16996
rect 42756 16940 42766 16996
rect 1810 16828 1820 16884
rect 1876 16828 5068 16884
rect 5124 16828 9660 16884
rect 9716 16828 11900 16884
rect 11956 16828 11966 16884
rect 13234 16828 13244 16884
rect 13300 16828 14588 16884
rect 14644 16828 14654 16884
rect 14812 16828 15820 16884
rect 15876 16828 17388 16884
rect 17444 16828 18060 16884
rect 18116 16828 18126 16884
rect 33506 16828 33516 16884
rect 33572 16828 34300 16884
rect 34356 16828 34366 16884
rect 47618 16828 47628 16884
rect 47684 16828 48748 16884
rect 48804 16828 48814 16884
rect 49410 16828 49420 16884
rect 49476 16828 50204 16884
rect 50260 16828 50270 16884
rect 18610 16716 18620 16772
rect 18676 16716 19628 16772
rect 19684 16716 19694 16772
rect 21522 16716 21532 16772
rect 21588 16716 22316 16772
rect 22372 16716 22382 16772
rect 23538 16716 23548 16772
rect 23604 16716 25564 16772
rect 25620 16716 25630 16772
rect 36418 16716 36428 16772
rect 36484 16716 36764 16772
rect 36820 16716 36830 16772
rect 50764 16716 50988 16772
rect 51044 16716 53228 16772
rect 53284 16716 53294 16772
rect 19628 16660 19684 16716
rect 50764 16660 50820 16716
rect 54200 16660 55000 16688
rect 17826 16604 17836 16660
rect 17892 16604 18508 16660
rect 18564 16604 18574 16660
rect 19628 16604 21644 16660
rect 21700 16604 22204 16660
rect 22260 16604 22652 16660
rect 22708 16604 23212 16660
rect 23268 16604 25900 16660
rect 25956 16604 25966 16660
rect 49970 16604 49980 16660
rect 50036 16604 50820 16660
rect 53106 16604 53116 16660
rect 53172 16604 55000 16660
rect 54200 16576 55000 16604
rect 6402 16492 6412 16548
rect 6468 16492 9884 16548
rect 9940 16492 9950 16548
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 38210 16380 38220 16436
rect 38276 16380 39452 16436
rect 39508 16380 39518 16436
rect 49074 16380 49084 16436
rect 49140 16380 49980 16436
rect 50036 16380 50046 16436
rect 12114 16268 12124 16324
rect 12180 16268 15036 16324
rect 15092 16268 16492 16324
rect 16548 16268 16558 16324
rect 34738 16268 34748 16324
rect 34804 16268 38668 16324
rect 38724 16268 38734 16324
rect 6514 16156 6524 16212
rect 6580 16156 7532 16212
rect 7588 16156 7598 16212
rect 16706 16156 16716 16212
rect 16772 16156 18172 16212
rect 18228 16156 20524 16212
rect 20580 16156 20590 16212
rect 29810 16156 29820 16212
rect 29876 16156 31948 16212
rect 38546 16156 38556 16212
rect 38612 16156 41020 16212
rect 41076 16156 42924 16212
rect 42980 16156 42990 16212
rect 43138 16156 43148 16212
rect 43204 16156 44828 16212
rect 44884 16156 44894 16212
rect 49942 16156 49980 16212
rect 50036 16156 50046 16212
rect 6178 16044 6188 16100
rect 6244 16044 7084 16100
rect 7140 16044 7308 16100
rect 7364 16044 7374 16100
rect 11778 16044 11788 16100
rect 11844 16044 12460 16100
rect 12516 16044 12526 16100
rect 16258 16044 16268 16100
rect 16324 16044 17500 16100
rect 17556 16044 17566 16100
rect 31892 15988 31948 16156
rect 36306 16044 36316 16100
rect 36372 16044 40796 16100
rect 40852 16044 40862 16100
rect 15586 15932 15596 15988
rect 15652 15932 17052 15988
rect 17108 15932 17388 15988
rect 17444 15932 17454 15988
rect 31892 15932 34860 15988
rect 34916 15932 36204 15988
rect 36260 15932 36270 15988
rect 38098 15932 38108 15988
rect 38164 15932 40684 15988
rect 40740 15932 40750 15988
rect 44482 15932 44492 15988
rect 44548 15932 46956 15988
rect 47012 15932 47022 15988
rect 11890 15820 11900 15876
rect 11956 15820 12684 15876
rect 12740 15820 15148 15876
rect 15204 15820 15214 15876
rect 35634 15820 35644 15876
rect 35700 15820 37772 15876
rect 37828 15820 37838 15876
rect 37986 15820 37996 15876
rect 38052 15820 41468 15876
rect 41524 15820 43932 15876
rect 43988 15820 43998 15876
rect 32396 15708 41468 15764
rect 41524 15708 43260 15764
rect 43316 15708 44044 15764
rect 44100 15708 44110 15764
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 32396 15540 32452 15708
rect 50546 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50830 15708
rect 38658 15596 38668 15652
rect 38724 15596 38734 15652
rect 42914 15596 42924 15652
rect 42980 15596 43484 15652
rect 43540 15596 43550 15652
rect 31378 15484 31388 15540
rect 31444 15484 32396 15540
rect 32452 15484 32462 15540
rect 38668 15428 38724 15596
rect 39526 15484 39564 15540
rect 39620 15484 39630 15540
rect 45826 15484 45836 15540
rect 45892 15484 46396 15540
rect 46452 15484 46462 15540
rect 47954 15484 47964 15540
rect 48020 15484 50204 15540
rect 50260 15484 50270 15540
rect 4946 15372 4956 15428
rect 5012 15372 7084 15428
rect 7140 15372 8316 15428
rect 8372 15372 8764 15428
rect 8820 15372 8830 15428
rect 13122 15372 13132 15428
rect 13188 15372 14364 15428
rect 14420 15372 14430 15428
rect 18610 15372 18620 15428
rect 18676 15372 19292 15428
rect 19348 15372 19740 15428
rect 19796 15372 19806 15428
rect 33964 15372 37100 15428
rect 37156 15372 38444 15428
rect 38500 15372 38510 15428
rect 38668 15372 39788 15428
rect 39844 15372 39854 15428
rect 42354 15372 42364 15428
rect 42420 15372 44604 15428
rect 44660 15372 44670 15428
rect 47058 15372 47068 15428
rect 47124 15372 47628 15428
rect 47684 15372 47694 15428
rect 2594 15260 2604 15316
rect 2660 15260 7532 15316
rect 7588 15260 7598 15316
rect 8082 15260 8092 15316
rect 8148 15260 8652 15316
rect 8708 15260 8718 15316
rect 9538 15260 9548 15316
rect 9604 15260 9884 15316
rect 9940 15260 9950 15316
rect 25330 15260 25340 15316
rect 25396 15260 25406 15316
rect 9426 15148 9436 15204
rect 9492 15148 9772 15204
rect 9828 15148 9838 15204
rect 14018 15148 14028 15204
rect 14084 15148 16492 15204
rect 16548 15148 16558 15204
rect 18722 15148 18732 15204
rect 18788 15148 18844 15204
rect 18900 15148 18910 15204
rect 25340 15092 25396 15260
rect 33964 15204 34020 15372
rect 34514 15260 34524 15316
rect 34580 15260 36988 15316
rect 37044 15260 37054 15316
rect 41234 15260 41244 15316
rect 41300 15260 42476 15316
rect 42532 15260 42812 15316
rect 42868 15260 43708 15316
rect 43764 15260 43774 15316
rect 50306 15260 50316 15316
rect 50372 15260 50988 15316
rect 51044 15260 51054 15316
rect 29250 15148 29260 15204
rect 29316 15148 33964 15204
rect 34020 15148 34030 15204
rect 34626 15148 34636 15204
rect 34692 15148 36540 15204
rect 36596 15148 36606 15204
rect 38322 15148 38332 15204
rect 38388 15148 43148 15204
rect 43204 15148 43428 15204
rect 43698 15148 43708 15204
rect 43764 15148 44380 15204
rect 44436 15148 44446 15204
rect 46396 15148 47068 15204
rect 47124 15148 47134 15204
rect 50428 15148 50652 15204
rect 50708 15148 50718 15204
rect 43372 15092 43428 15148
rect 46396 15092 46452 15148
rect 50428 15092 50484 15148
rect 10434 15036 10444 15092
rect 10500 15036 11116 15092
rect 11172 15036 15148 15092
rect 16482 15036 16492 15092
rect 16548 15036 16828 15092
rect 16884 15036 24108 15092
rect 24164 15036 25396 15092
rect 30930 15036 30940 15092
rect 30996 15036 31612 15092
rect 31668 15036 32172 15092
rect 32228 15036 32238 15092
rect 43362 15036 43372 15092
rect 43428 15036 43438 15092
rect 43670 15036 43708 15092
rect 43764 15036 43774 15092
rect 46386 15036 46396 15092
rect 46452 15036 46462 15092
rect 49074 15036 49084 15092
rect 49140 15036 50484 15092
rect 15092 14980 15148 15036
rect 15092 14924 16604 14980
rect 16660 14924 16670 14980
rect 38770 14924 38780 14980
rect 38836 14924 39900 14980
rect 39956 14924 39966 14980
rect 40226 14924 40236 14980
rect 40292 14924 46060 14980
rect 46116 14924 46126 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 32498 14700 32508 14756
rect 32564 14700 33068 14756
rect 33124 14700 33628 14756
rect 33684 14700 33694 14756
rect 38882 14588 38892 14644
rect 38948 14588 40684 14644
rect 40740 14588 40750 14644
rect 49970 14588 49980 14644
rect 50036 14588 52668 14644
rect 52724 14588 52734 14644
rect 11330 14476 11340 14532
rect 11396 14476 12012 14532
rect 12068 14476 12078 14532
rect 16594 14476 16604 14532
rect 16660 14476 17276 14532
rect 17332 14476 17342 14532
rect 18386 14476 18396 14532
rect 18452 14476 19068 14532
rect 19124 14476 20636 14532
rect 20692 14476 20702 14532
rect 34402 14476 34412 14532
rect 34468 14476 35868 14532
rect 35924 14476 35934 14532
rect 48850 14476 48860 14532
rect 48916 14476 49644 14532
rect 49700 14476 49710 14532
rect 31266 14364 31276 14420
rect 31332 14364 32284 14420
rect 32340 14364 32350 14420
rect 33170 14364 33180 14420
rect 33236 14364 35308 14420
rect 35364 14364 35374 14420
rect 38098 14364 38108 14420
rect 38164 14364 41916 14420
rect 41972 14364 42588 14420
rect 42644 14364 42654 14420
rect 45714 14364 45724 14420
rect 45780 14364 46508 14420
rect 46564 14364 46574 14420
rect 6178 14252 6188 14308
rect 6244 14252 7084 14308
rect 7140 14252 7150 14308
rect 8082 14252 8092 14308
rect 8148 14252 10220 14308
rect 10276 14252 12124 14308
rect 12180 14252 12190 14308
rect 16930 14252 16940 14308
rect 16996 14252 17164 14308
rect 17220 14252 18844 14308
rect 18900 14252 18910 14308
rect 26114 14252 26124 14308
rect 26180 14252 26572 14308
rect 26628 14252 26908 14308
rect 27906 14252 27916 14308
rect 27972 14252 31388 14308
rect 31444 14252 31454 14308
rect 32162 14252 32172 14308
rect 32228 14252 33068 14308
rect 33124 14252 33134 14308
rect 39666 14252 39676 14308
rect 39732 14252 40796 14308
rect 40852 14252 40862 14308
rect 41234 14252 41244 14308
rect 41300 14252 42252 14308
rect 42308 14252 46172 14308
rect 46228 14252 46238 14308
rect 46386 14252 46396 14308
rect 46452 14252 46844 14308
rect 46900 14252 46910 14308
rect 49074 14252 49084 14308
rect 49140 14252 50092 14308
rect 50148 14252 50158 14308
rect 26852 14196 26908 14252
rect 46396 14196 46452 14252
rect 26852 14140 31948 14196
rect 32386 14140 32396 14196
rect 32452 14140 40012 14196
rect 40068 14140 41916 14196
rect 41972 14140 41982 14196
rect 46050 14140 46060 14196
rect 46116 14140 46452 14196
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 31892 14084 31948 14140
rect 46060 14084 46116 14140
rect 50546 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50830 14140
rect 31892 14028 46116 14084
rect 54200 13972 55000 14000
rect 6402 13916 6412 13972
rect 6468 13916 7308 13972
rect 7364 13916 11004 13972
rect 11060 13916 11070 13972
rect 16146 13916 16156 13972
rect 16212 13916 17724 13972
rect 17780 13916 26908 13972
rect 32498 13916 32508 13972
rect 32564 13916 32956 13972
rect 33012 13916 33852 13972
rect 33908 13916 33918 13972
rect 46134 13916 46172 13972
rect 46228 13916 46238 13972
rect 52210 13916 52220 13972
rect 52276 13916 53228 13972
rect 53284 13916 55000 13972
rect 26852 13860 26908 13916
rect 54200 13888 55000 13916
rect 16370 13804 16380 13860
rect 16436 13804 17052 13860
rect 17108 13804 17612 13860
rect 17668 13804 18284 13860
rect 18340 13804 18350 13860
rect 26852 13804 31164 13860
rect 31220 13804 31230 13860
rect 31826 13804 31836 13860
rect 31892 13804 33180 13860
rect 33236 13804 33246 13860
rect 11666 13692 11676 13748
rect 11732 13692 12348 13748
rect 12404 13692 12414 13748
rect 14354 13692 14364 13748
rect 14420 13692 15932 13748
rect 15988 13692 15998 13748
rect 18498 13692 18508 13748
rect 18564 13692 20300 13748
rect 20356 13692 27692 13748
rect 27748 13692 27758 13748
rect 31938 13692 31948 13748
rect 32004 13692 32014 13748
rect 15932 13636 15988 13692
rect 2482 13580 2492 13636
rect 2548 13580 6076 13636
rect 6132 13580 6142 13636
rect 15932 13580 18732 13636
rect 18788 13580 18798 13636
rect 19058 13580 19068 13636
rect 19124 13580 19516 13636
rect 19572 13580 19582 13636
rect 25330 13580 25340 13636
rect 25396 13580 26460 13636
rect 26516 13580 26796 13636
rect 26852 13580 26862 13636
rect 7186 13468 7196 13524
rect 7252 13468 8092 13524
rect 8148 13468 8158 13524
rect 10658 13468 10668 13524
rect 10724 13468 11564 13524
rect 11620 13468 11630 13524
rect 18834 13468 18844 13524
rect 18900 13468 19404 13524
rect 19460 13468 19470 13524
rect 21858 13468 21868 13524
rect 21924 13468 22876 13524
rect 22932 13468 22942 13524
rect 14466 13356 14476 13412
rect 14532 13356 14812 13412
rect 14868 13356 15484 13412
rect 15540 13356 15550 13412
rect 25218 13356 25228 13412
rect 25284 13356 26348 13412
rect 26404 13356 26414 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 4834 13244 4844 13300
rect 4900 13244 6412 13300
rect 6468 13244 6478 13300
rect 26852 13244 31052 13300
rect 31108 13244 31118 13300
rect 6178 13132 6188 13188
rect 6244 13132 8316 13188
rect 8372 13132 8382 13188
rect 7196 13076 7252 13132
rect 4946 13020 4956 13076
rect 5012 13020 5740 13076
rect 5796 13020 5806 13076
rect 7186 13020 7196 13076
rect 7252 13020 7262 13076
rect 10994 13020 11004 13076
rect 11060 13020 11900 13076
rect 11956 13020 26684 13076
rect 26740 13020 26750 13076
rect 26852 12964 26908 13244
rect 31948 13188 32004 13692
rect 49634 13580 49644 13636
rect 49700 13580 53228 13636
rect 53284 13580 53294 13636
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 39218 13244 39228 13300
rect 39284 13244 40460 13300
rect 40516 13244 40526 13300
rect 46834 13244 46844 13300
rect 46900 13244 47404 13300
rect 47460 13244 48636 13300
rect 48692 13244 48702 13300
rect 31948 13132 35644 13188
rect 35700 13132 38108 13188
rect 38164 13132 38174 13188
rect 27682 13020 27692 13076
rect 27748 13020 28588 13076
rect 28644 13020 28654 13076
rect 5058 12908 5068 12964
rect 5124 12908 5964 12964
rect 6020 12908 6860 12964
rect 6916 12908 6926 12964
rect 12114 12908 12124 12964
rect 12180 12908 13916 12964
rect 13972 12908 13982 12964
rect 14242 12908 14252 12964
rect 14308 12908 15148 12964
rect 15204 12908 26908 12964
rect 38322 12908 38332 12964
rect 38388 12908 40012 12964
rect 40068 12908 40078 12964
rect 42242 12908 42252 12964
rect 42308 12908 43148 12964
rect 43204 12908 43708 12964
rect 43764 12908 43774 12964
rect 4946 12796 4956 12852
rect 5012 12796 5628 12852
rect 5684 12796 5694 12852
rect 22418 12796 22428 12852
rect 22484 12796 23996 12852
rect 24052 12796 24062 12852
rect 5926 12684 5964 12740
rect 6020 12684 6030 12740
rect 33058 12684 33068 12740
rect 33124 12684 35532 12740
rect 35588 12684 35868 12740
rect 35924 12684 35934 12740
rect 36082 12684 36092 12740
rect 36148 12684 37772 12740
rect 37828 12684 38556 12740
rect 38612 12684 38622 12740
rect 39750 12684 39788 12740
rect 39844 12684 39854 12740
rect 45602 12684 45612 12740
rect 45668 12684 46284 12740
rect 46340 12684 46350 12740
rect 48972 12684 50764 12740
rect 50820 12684 50830 12740
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 48972 12516 49028 12684
rect 50546 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50830 12572
rect 38612 12460 45388 12516
rect 45444 12460 45724 12516
rect 45780 12460 45790 12516
rect 48962 12460 48972 12516
rect 49028 12460 49038 12516
rect 38612 12404 38668 12460
rect 15092 12348 25228 12404
rect 25284 12348 25294 12404
rect 25526 12348 25564 12404
rect 25620 12348 25630 12404
rect 27122 12348 27132 12404
rect 27188 12348 28812 12404
rect 28868 12348 29260 12404
rect 29316 12348 29326 12404
rect 34962 12348 34972 12404
rect 35028 12348 38668 12404
rect 40338 12348 40348 12404
rect 40404 12348 41020 12404
rect 41076 12348 41580 12404
rect 41636 12348 41646 12404
rect 5842 12236 5852 12292
rect 5908 12236 9548 12292
rect 9604 12236 9614 12292
rect 14130 12236 14140 12292
rect 14196 12236 14812 12292
rect 14868 12236 14878 12292
rect 15092 12180 15148 12348
rect 40348 12180 40404 12348
rect 46946 12236 46956 12292
rect 47012 12236 52444 12292
rect 52500 12236 52510 12292
rect 9202 12124 9212 12180
rect 9268 12124 10108 12180
rect 10164 12124 10174 12180
rect 12450 12124 12460 12180
rect 12516 12124 13468 12180
rect 13524 12124 15148 12180
rect 20738 12124 20748 12180
rect 20804 12124 21868 12180
rect 21924 12124 21934 12180
rect 22306 12124 22316 12180
rect 22372 12124 23884 12180
rect 23940 12124 23950 12180
rect 24210 12124 24220 12180
rect 24276 12124 25116 12180
rect 25172 12124 27244 12180
rect 27300 12124 27310 12180
rect 35970 12124 35980 12180
rect 36036 12124 37100 12180
rect 37156 12124 40404 12180
rect 1810 12012 1820 12068
rect 1876 12012 4844 12068
rect 4900 12012 4910 12068
rect 12898 12012 12908 12068
rect 12964 12012 14476 12068
rect 14532 12012 14542 12068
rect 35186 12012 35196 12068
rect 35252 12012 36428 12068
rect 36484 12012 36494 12068
rect 8306 11900 8316 11956
rect 8372 11900 10332 11956
rect 10388 11900 12572 11956
rect 12628 11900 12638 11956
rect 15250 11900 15260 11956
rect 15316 11900 19180 11956
rect 19236 11900 19246 11956
rect 33954 11900 33964 11956
rect 34020 11900 35420 11956
rect 35476 11900 35486 11956
rect 36530 11788 36540 11844
rect 36596 11788 38220 11844
rect 38276 11788 45948 11844
rect 46004 11788 48972 11844
rect 49028 11788 49038 11844
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 13346 11676 13356 11732
rect 13412 11676 14588 11732
rect 14644 11676 14654 11732
rect 21410 11676 21420 11732
rect 21476 11676 22204 11732
rect 22260 11676 22270 11732
rect 44818 11676 44828 11732
rect 44884 11676 46172 11732
rect 46228 11676 46620 11732
rect 46676 11676 46686 11732
rect 14354 11564 14364 11620
rect 14420 11564 15932 11620
rect 15988 11564 15998 11620
rect 5954 11452 5964 11508
rect 6020 11452 7868 11508
rect 7924 11452 8204 11508
rect 8260 11452 8270 11508
rect 15138 11452 15148 11508
rect 15204 11452 16604 11508
rect 16660 11452 16670 11508
rect 29922 11452 29932 11508
rect 29988 11452 31836 11508
rect 31892 11452 31902 11508
rect 6626 11340 6636 11396
rect 6692 11340 9380 11396
rect 14802 11340 14812 11396
rect 14868 11340 15820 11396
rect 15876 11340 18844 11396
rect 18900 11340 18910 11396
rect 40786 11340 40796 11396
rect 40852 11340 41916 11396
rect 41972 11340 41982 11396
rect 9324 11284 9380 11340
rect 54200 11284 55000 11312
rect 4274 11228 4284 11284
rect 4340 11228 8652 11284
rect 8708 11228 8718 11284
rect 9314 11228 9324 11284
rect 9380 11228 10892 11284
rect 10948 11228 10958 11284
rect 11666 11228 11676 11284
rect 11732 11228 12796 11284
rect 12852 11228 14028 11284
rect 14084 11228 15148 11284
rect 15204 11228 15214 11284
rect 26226 11228 26236 11284
rect 26292 11228 26684 11284
rect 26740 11228 28028 11284
rect 28084 11228 31500 11284
rect 31556 11228 32732 11284
rect 32788 11228 32798 11284
rect 45350 11228 45388 11284
rect 45444 11228 45454 11284
rect 45574 11228 45612 11284
rect 45668 11228 45678 11284
rect 53218 11228 53228 11284
rect 53284 11228 55000 11284
rect 54200 11200 55000 11228
rect 2482 11116 2492 11172
rect 2548 11116 5740 11172
rect 5796 11116 5806 11172
rect 6066 11116 6076 11172
rect 6132 11116 6972 11172
rect 7028 11116 7038 11172
rect 14354 11116 14364 11172
rect 14420 11116 15260 11172
rect 15316 11116 15326 11172
rect 21522 11116 21532 11172
rect 21588 11116 24780 11172
rect 24836 11116 25340 11172
rect 25396 11116 25406 11172
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 50546 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50830 11004
rect 10994 10892 11004 10948
rect 11060 10892 12124 10948
rect 12180 10892 13300 10948
rect 27346 10892 27356 10948
rect 27412 10892 27916 10948
rect 27972 10892 29820 10948
rect 29876 10892 37436 10948
rect 37492 10892 37502 10948
rect 44146 10892 44156 10948
rect 44212 10892 45052 10948
rect 45108 10892 45118 10948
rect 13244 10836 13300 10892
rect 4162 10780 4172 10836
rect 4228 10780 4620 10836
rect 4676 10780 5068 10836
rect 5124 10780 5134 10836
rect 7746 10780 7756 10836
rect 7812 10780 10892 10836
rect 10948 10780 10958 10836
rect 12002 10780 12012 10836
rect 12068 10780 12078 10836
rect 13234 10780 13244 10836
rect 13300 10780 19068 10836
rect 19124 10780 19134 10836
rect 12012 10724 12068 10780
rect 10658 10668 10668 10724
rect 10724 10668 12068 10724
rect 12562 10556 12572 10612
rect 12628 10556 13916 10612
rect 13972 10556 13982 10612
rect 45042 10556 45052 10612
rect 45108 10556 45724 10612
rect 45780 10556 46396 10612
rect 46452 10556 46462 10612
rect 46722 10556 46732 10612
rect 46788 10556 47180 10612
rect 47236 10556 49196 10612
rect 49252 10556 49262 10612
rect 11442 10444 11452 10500
rect 11508 10444 13356 10500
rect 13412 10444 13422 10500
rect 36194 10332 36204 10388
rect 36260 10332 42700 10388
rect 42756 10332 42766 10388
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 7186 10108 7196 10164
rect 7252 10108 8428 10164
rect 31490 10108 31500 10164
rect 31556 10108 34972 10164
rect 35028 10108 35038 10164
rect 41682 10108 41692 10164
rect 41748 10108 44492 10164
rect 44548 10108 45500 10164
rect 45556 10108 45566 10164
rect 8372 10052 8428 10108
rect 8372 9996 30268 10052
rect 30324 9996 30334 10052
rect 34850 9996 34860 10052
rect 34916 9996 35868 10052
rect 35924 9996 37660 10052
rect 37716 9996 37726 10052
rect 41010 9996 41020 10052
rect 41076 9996 41916 10052
rect 41972 9996 41982 10052
rect 46162 9996 46172 10052
rect 46228 9996 52892 10052
rect 52948 9996 52958 10052
rect 21298 9884 21308 9940
rect 21364 9884 22092 9940
rect 22148 9884 22764 9940
rect 22820 9884 25116 9940
rect 25172 9884 25182 9940
rect 25778 9884 25788 9940
rect 25844 9884 26460 9940
rect 26516 9884 42700 9940
rect 42756 9884 42766 9940
rect 49298 9884 49308 9940
rect 49364 9884 50764 9940
rect 50820 9884 50830 9940
rect 4162 9772 4172 9828
rect 4228 9772 6972 9828
rect 7028 9772 7644 9828
rect 7700 9772 7710 9828
rect 32498 9772 32508 9828
rect 32564 9772 33852 9828
rect 33908 9772 35308 9828
rect 35364 9772 35374 9828
rect 38210 9772 38220 9828
rect 38276 9772 38668 9828
rect 38724 9772 39676 9828
rect 39732 9772 39742 9828
rect 44258 9772 44268 9828
rect 44324 9772 45052 9828
rect 45108 9772 45118 9828
rect 45378 9772 45388 9828
rect 45444 9772 48860 9828
rect 48916 9772 49420 9828
rect 49476 9772 49486 9828
rect 32946 9660 32956 9716
rect 33012 9660 33516 9716
rect 33572 9660 33582 9716
rect 35970 9660 35980 9716
rect 36036 9660 39900 9716
rect 39956 9660 39966 9716
rect 43586 9660 43596 9716
rect 43652 9660 47964 9716
rect 48020 9660 48030 9716
rect 49186 9660 49196 9716
rect 49252 9660 49868 9716
rect 49924 9660 53340 9716
rect 53396 9660 53406 9716
rect 47964 9604 48020 9660
rect 13682 9548 13692 9604
rect 13748 9548 15484 9604
rect 15540 9548 16716 9604
rect 16772 9548 16782 9604
rect 37090 9548 37100 9604
rect 37156 9548 37660 9604
rect 37716 9548 39228 9604
rect 39284 9548 39294 9604
rect 42690 9548 42700 9604
rect 42756 9548 44268 9604
rect 44324 9548 45164 9604
rect 45220 9548 45230 9604
rect 46610 9548 46620 9604
rect 46676 9548 46956 9604
rect 47012 9548 47022 9604
rect 47964 9548 49532 9604
rect 49588 9548 49598 9604
rect 37100 9492 37156 9548
rect 31154 9436 31164 9492
rect 31220 9436 37156 9492
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 50546 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50830 9436
rect 7746 9212 7756 9268
rect 7812 9212 9884 9268
rect 9940 9212 11340 9268
rect 11396 9212 11406 9268
rect 35634 9212 35644 9268
rect 35700 9212 37996 9268
rect 38052 9212 38062 9268
rect 46162 9212 46172 9268
rect 46228 9212 48524 9268
rect 48580 9212 48590 9268
rect 39890 9100 39900 9156
rect 39956 9100 41244 9156
rect 41300 9100 41916 9156
rect 41972 9100 41982 9156
rect 43362 9100 43372 9156
rect 43428 9100 46620 9156
rect 46676 9100 46686 9156
rect 31892 8988 40124 9044
rect 40180 8988 40190 9044
rect 41458 8988 41468 9044
rect 41524 8988 45052 9044
rect 45108 8988 45388 9044
rect 45444 8988 45454 9044
rect 20290 8876 20300 8932
rect 20356 8876 22204 8932
rect 22260 8876 22270 8932
rect 29362 8876 29372 8932
rect 29428 8876 30716 8932
rect 30772 8876 30782 8932
rect 31892 8820 31948 8988
rect 33394 8876 33404 8932
rect 33460 8876 35532 8932
rect 35588 8876 35598 8932
rect 42802 8876 42812 8932
rect 42868 8876 44380 8932
rect 44436 8876 44446 8932
rect 30594 8764 30604 8820
rect 30660 8764 31948 8820
rect 45574 8652 45612 8708
rect 45668 8652 45678 8708
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 54200 8596 55000 8624
rect 42242 8540 42252 8596
rect 42308 8540 43372 8596
rect 43428 8540 43438 8596
rect 53218 8540 53228 8596
rect 53284 8540 55000 8596
rect 54200 8512 55000 8540
rect 11330 8428 11340 8484
rect 11396 8428 13356 8484
rect 13412 8428 16828 8484
rect 16884 8428 16894 8484
rect 20178 8428 20188 8484
rect 20244 8428 20972 8484
rect 21028 8428 21038 8484
rect 26348 8428 26572 8484
rect 26628 8428 27020 8484
rect 27076 8428 31276 8484
rect 31332 8428 31342 8484
rect 40338 8428 40348 8484
rect 40404 8428 43036 8484
rect 43092 8428 45612 8484
rect 45668 8428 45678 8484
rect 18162 8316 18172 8372
rect 18228 8316 19404 8372
rect 19460 8316 19470 8372
rect 7858 8204 7868 8260
rect 7924 8204 8988 8260
rect 9044 8204 9054 8260
rect 19618 8204 19628 8260
rect 19684 8204 20524 8260
rect 20580 8204 21980 8260
rect 22036 8204 22046 8260
rect 22642 8204 22652 8260
rect 22708 8204 25564 8260
rect 25620 8204 25900 8260
rect 25956 8204 25966 8260
rect 7298 8092 7308 8148
rect 7364 8092 8876 8148
rect 8932 8092 8942 8148
rect 19730 8092 19740 8148
rect 19796 8092 20412 8148
rect 20468 8092 20478 8148
rect 26348 8036 26404 8428
rect 44818 8316 44828 8372
rect 44884 8316 45276 8372
rect 45332 8316 46844 8372
rect 46900 8316 48636 8372
rect 48692 8316 48702 8372
rect 37314 8204 37324 8260
rect 37380 8204 47740 8260
rect 47796 8204 49084 8260
rect 49140 8204 49150 8260
rect 49644 8092 50540 8148
rect 50596 8092 50606 8148
rect 49644 8036 49700 8092
rect 8082 7980 8092 8036
rect 8148 7980 9548 8036
rect 9604 7980 10780 8036
rect 10836 7980 10846 8036
rect 20738 7980 20748 8036
rect 20804 7980 22092 8036
rect 22148 7980 22158 8036
rect 23090 7980 23100 8036
rect 23156 7980 24780 8036
rect 24836 7980 26348 8036
rect 26404 7980 26414 8036
rect 26852 7980 29036 8036
rect 29092 7980 29102 8036
rect 37986 7980 37996 8036
rect 38052 7980 39564 8036
rect 39620 7980 39630 8036
rect 45378 7980 45388 8036
rect 45444 7980 48188 8036
rect 48244 7980 48524 8036
rect 48580 7980 48590 8036
rect 49634 7980 49644 8036
rect 49700 7980 49710 8036
rect 50372 7980 52668 8036
rect 52724 7980 52734 8036
rect 26852 7924 26908 7980
rect 20290 7868 20300 7924
rect 20356 7868 22428 7924
rect 22484 7868 26908 7924
rect 41794 7868 41804 7924
rect 41860 7868 42476 7924
rect 42532 7868 46060 7924
rect 46116 7868 46126 7924
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 50372 7812 50428 7980
rect 50546 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50830 7868
rect 38322 7756 38332 7812
rect 38388 7756 47068 7812
rect 47124 7756 47134 7812
rect 49410 7756 49420 7812
rect 49476 7756 50428 7812
rect 8306 7644 8316 7700
rect 8372 7644 8988 7700
rect 9044 7644 9054 7700
rect 19506 7644 19516 7700
rect 19572 7644 20860 7700
rect 20916 7644 23548 7700
rect 23604 7644 23614 7700
rect 29698 7644 29708 7700
rect 29764 7644 30268 7700
rect 30324 7644 31948 7700
rect 32274 7644 32284 7700
rect 32340 7644 33180 7700
rect 33236 7644 40852 7700
rect 44034 7644 44044 7700
rect 44100 7644 45500 7700
rect 45556 7644 45566 7700
rect 31892 7588 31948 7644
rect 12114 7532 12124 7588
rect 12180 7532 14140 7588
rect 14196 7532 14206 7588
rect 18274 7532 18284 7588
rect 18340 7532 19628 7588
rect 19684 7532 19694 7588
rect 25666 7532 25676 7588
rect 25732 7532 27580 7588
rect 27636 7532 30324 7588
rect 31892 7532 37548 7588
rect 37604 7532 37614 7588
rect 30268 7476 30324 7532
rect 40796 7476 40852 7644
rect 47954 7532 47964 7588
rect 48020 7532 49532 7588
rect 49588 7532 49598 7588
rect 19506 7420 19516 7476
rect 19572 7420 19852 7476
rect 19908 7420 20300 7476
rect 20356 7420 20366 7476
rect 22306 7420 22316 7476
rect 22372 7420 30044 7476
rect 30100 7420 30110 7476
rect 30268 7420 35756 7476
rect 35812 7420 35822 7476
rect 40786 7420 40796 7476
rect 40852 7420 40862 7476
rect 45154 7420 45164 7476
rect 45220 7420 46284 7476
rect 46340 7420 46350 7476
rect 48178 7420 48188 7476
rect 48244 7420 49308 7476
rect 49364 7420 49374 7476
rect 19954 7308 19964 7364
rect 20020 7308 20636 7364
rect 20692 7308 20702 7364
rect 38770 7308 38780 7364
rect 38836 7308 44044 7364
rect 44100 7308 44110 7364
rect 23538 7084 23548 7140
rect 23604 7084 25788 7140
rect 25844 7084 26908 7140
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 26852 6916 26908 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 48738 6972 48748 7028
rect 48804 6972 49308 7028
rect 49364 6972 49374 7028
rect 26852 6860 33292 6916
rect 33348 6860 33358 6916
rect 48962 6860 48972 6916
rect 49028 6860 49868 6916
rect 49924 6860 49934 6916
rect 16146 6748 16156 6804
rect 16212 6748 20748 6804
rect 20804 6748 20814 6804
rect 32162 6748 32172 6804
rect 32228 6748 36204 6804
rect 36260 6748 36270 6804
rect 42476 6748 45388 6804
rect 45444 6748 45454 6804
rect 47730 6748 47740 6804
rect 47796 6748 48188 6804
rect 48244 6748 49084 6804
rect 49140 6748 50316 6804
rect 50372 6748 50382 6804
rect 42476 6692 42532 6748
rect 13570 6636 13580 6692
rect 13636 6636 14700 6692
rect 14756 6636 15036 6692
rect 15092 6636 15372 6692
rect 15428 6636 15438 6692
rect 38210 6636 38220 6692
rect 38276 6636 38780 6692
rect 38836 6636 38846 6692
rect 42466 6636 42476 6692
rect 42532 6636 42542 6692
rect 48402 6636 48412 6692
rect 48468 6636 49644 6692
rect 49700 6636 49710 6692
rect 32498 6524 32508 6580
rect 32564 6524 33628 6580
rect 33684 6524 33694 6580
rect 37426 6524 37436 6580
rect 37492 6524 38332 6580
rect 38388 6524 39228 6580
rect 39284 6524 39294 6580
rect 41794 6524 41804 6580
rect 41860 6524 42028 6580
rect 42084 6524 45164 6580
rect 45220 6524 45230 6580
rect 45490 6524 45500 6580
rect 45556 6524 46620 6580
rect 46676 6524 47404 6580
rect 47460 6524 47470 6580
rect 50372 6524 52668 6580
rect 52724 6524 52734 6580
rect 50372 6468 50428 6524
rect 21634 6412 21644 6468
rect 21700 6412 22876 6468
rect 22932 6412 24444 6468
rect 24500 6412 26796 6468
rect 26852 6412 26862 6468
rect 46050 6412 46060 6468
rect 46116 6412 46732 6468
rect 46788 6412 50428 6468
rect 51314 6412 51324 6468
rect 51380 6412 51996 6468
rect 52052 6412 52062 6468
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 50546 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50830 6300
rect 22418 6188 22428 6244
rect 22484 6188 27580 6244
rect 27636 6188 27646 6244
rect 19506 6076 19516 6132
rect 19572 6076 19740 6132
rect 19796 6076 19806 6132
rect 20178 6076 20188 6132
rect 20244 6076 21756 6132
rect 21812 6076 21822 6132
rect 27458 6076 27468 6132
rect 27524 6076 31724 6132
rect 31780 6076 33068 6132
rect 33124 6076 33134 6132
rect 41682 6076 41692 6132
rect 41748 6076 42364 6132
rect 42420 6076 42430 6132
rect 44930 6076 44940 6132
rect 44996 6076 51548 6132
rect 51604 6076 51614 6132
rect 19954 5964 19964 6020
rect 20020 5964 20300 6020
rect 20356 5964 21308 6020
rect 21364 5964 21374 6020
rect 54200 5908 55000 5936
rect 17378 5852 17388 5908
rect 17444 5852 19628 5908
rect 19684 5852 19694 5908
rect 21410 5852 21420 5908
rect 21476 5852 22652 5908
rect 22708 5852 28140 5908
rect 28196 5852 29260 5908
rect 29316 5852 29708 5908
rect 29764 5852 29774 5908
rect 33730 5852 33740 5908
rect 33796 5852 35980 5908
rect 36036 5852 36046 5908
rect 36194 5852 36204 5908
rect 36260 5852 37212 5908
rect 37268 5852 43260 5908
rect 43316 5852 43326 5908
rect 51986 5852 51996 5908
rect 52052 5852 55000 5908
rect 54200 5824 55000 5852
rect 50372 5740 51100 5796
rect 51156 5740 51166 5796
rect 50372 5684 50428 5740
rect 15250 5628 15260 5684
rect 15316 5628 18844 5684
rect 18900 5628 18910 5684
rect 49970 5628 49980 5684
rect 50036 5628 50428 5684
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19170 5292 19180 5348
rect 19236 5292 21532 5348
rect 21588 5292 21598 5348
rect 30146 5292 30156 5348
rect 30212 5292 31500 5348
rect 31556 5292 31566 5348
rect 29586 5180 29596 5236
rect 29652 5180 30380 5236
rect 30436 5180 30446 5236
rect 32946 5180 32956 5236
rect 33012 5180 36428 5236
rect 36484 5180 36876 5236
rect 36932 5180 36942 5236
rect 14690 5068 14700 5124
rect 14756 5068 16828 5124
rect 16884 5068 17836 5124
rect 17892 5068 17902 5124
rect 18946 5068 18956 5124
rect 19012 5068 22540 5124
rect 22596 5068 25228 5124
rect 25284 5068 25788 5124
rect 25844 5068 25854 5124
rect 26114 5068 26124 5124
rect 26180 5068 28252 5124
rect 28308 5068 28318 5124
rect 42130 5068 42140 5124
rect 42196 5068 43820 5124
rect 43876 5068 46284 5124
rect 46340 5068 46350 5124
rect 46498 5068 46508 5124
rect 46564 5068 48636 5124
rect 48692 5068 53228 5124
rect 53284 5068 53294 5124
rect 28354 4956 28364 5012
rect 28420 4956 31612 5012
rect 31668 4956 32172 5012
rect 32228 4956 32238 5012
rect 44034 4956 44044 5012
rect 44100 4956 52668 5012
rect 52724 4956 52734 5012
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 50546 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50830 4732
rect 31892 4620 37100 4676
rect 37156 4620 37166 4676
rect 31892 4452 31948 4620
rect 36978 4508 36988 4564
rect 37044 4508 40236 4564
rect 40292 4508 40572 4564
rect 40628 4508 41020 4564
rect 41076 4508 41086 4564
rect 14354 4396 14364 4452
rect 14420 4396 14924 4452
rect 14980 4396 31948 4452
rect 33170 4396 33180 4452
rect 33236 4396 33852 4452
rect 33908 4396 33918 4452
rect 48178 4396 48188 4452
rect 48244 4396 50876 4452
rect 50932 4396 50942 4452
rect 21634 4284 21644 4340
rect 21700 4284 24668 4340
rect 24724 4284 25228 4340
rect 25284 4284 26348 4340
rect 26404 4284 29260 4340
rect 29316 4284 29326 4340
rect 44258 4284 44268 4340
rect 44324 4284 47516 4340
rect 47572 4284 49084 4340
rect 49140 4284 50316 4340
rect 50372 4284 51660 4340
rect 51716 4284 51726 4340
rect 3714 4172 3724 4228
rect 3780 4172 28812 4228
rect 28868 4172 28878 4228
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 31892 3724 38892 3780
rect 38948 3724 39788 3780
rect 39844 3724 39854 3780
rect 31892 3668 31948 3724
rect 11890 3612 11900 3668
rect 11956 3612 12460 3668
rect 12516 3612 31948 3668
rect 34066 3612 34076 3668
rect 34132 3612 36988 3668
rect 37044 3612 37054 3668
rect 50418 3612 50428 3668
rect 50484 3612 51996 3668
rect 52052 3612 52062 3668
rect 10770 3500 10780 3556
rect 10836 3500 35532 3556
rect 35588 3500 35980 3556
rect 36036 3500 36046 3556
rect 46946 3500 46956 3556
rect 47012 3500 47628 3556
rect 47684 3500 47694 3556
rect 7186 3388 7196 3444
rect 7252 3388 10108 3444
rect 10164 3388 10174 3444
rect 38546 3388 38556 3444
rect 38612 3388 39340 3444
rect 39396 3388 39788 3444
rect 39844 3388 39854 3444
rect 45378 3388 45388 3444
rect 45444 3388 47460 3444
rect 47404 3332 47460 3388
rect 16146 3276 16156 3332
rect 16212 3276 16940 3332
rect 16996 3276 17006 3332
rect 47394 3276 47404 3332
rect 47460 3276 47470 3332
rect 54200 3220 55000 3248
rect 52434 3164 52444 3220
rect 52500 3164 53228 3220
rect 53284 3164 55000 3220
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
rect 50546 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50830 3164
rect 54200 3136 55000 3164
<< via3 >>
rect 19836 51716 19892 51772
rect 19940 51716 19996 51772
rect 20044 51716 20100 51772
rect 50556 51716 50612 51772
rect 50660 51716 50716 51772
rect 50764 51716 50820 51772
rect 4476 50932 4532 50988
rect 4580 50932 4636 50988
rect 4684 50932 4740 50988
rect 35196 50932 35252 50988
rect 35300 50932 35356 50988
rect 35404 50932 35460 50988
rect 19836 50148 19892 50204
rect 19940 50148 19996 50204
rect 20044 50148 20100 50204
rect 50556 50148 50612 50204
rect 50660 50148 50716 50204
rect 50764 50148 50820 50204
rect 4476 49364 4532 49420
rect 4580 49364 4636 49420
rect 4684 49364 4740 49420
rect 35196 49364 35252 49420
rect 35300 49364 35356 49420
rect 35404 49364 35460 49420
rect 19836 48580 19892 48636
rect 19940 48580 19996 48636
rect 20044 48580 20100 48636
rect 50556 48580 50612 48636
rect 50660 48580 50716 48636
rect 50764 48580 50820 48636
rect 4476 47796 4532 47852
rect 4580 47796 4636 47852
rect 4684 47796 4740 47852
rect 35196 47796 35252 47852
rect 35300 47796 35356 47852
rect 35404 47796 35460 47852
rect 19836 47012 19892 47068
rect 19940 47012 19996 47068
rect 20044 47012 20100 47068
rect 50556 47012 50612 47068
rect 50660 47012 50716 47068
rect 50764 47012 50820 47068
rect 47068 46620 47124 46676
rect 4476 46228 4532 46284
rect 4580 46228 4636 46284
rect 4684 46228 4740 46284
rect 35196 46228 35252 46284
rect 35300 46228 35356 46284
rect 35404 46228 35460 46284
rect 19180 46172 19236 46228
rect 19836 45444 19892 45500
rect 19940 45444 19996 45500
rect 20044 45444 20100 45500
rect 50556 45444 50612 45500
rect 50660 45444 50716 45500
rect 50764 45444 50820 45500
rect 19068 45164 19124 45220
rect 4476 44660 4532 44716
rect 4580 44660 4636 44716
rect 4684 44660 4740 44716
rect 35196 44660 35252 44716
rect 35300 44660 35356 44716
rect 35404 44660 35460 44716
rect 19836 43876 19892 43932
rect 19940 43876 19996 43932
rect 20044 43876 20100 43932
rect 50556 43876 50612 43932
rect 50660 43876 50716 43932
rect 50764 43876 50820 43932
rect 4476 43092 4532 43148
rect 4580 43092 4636 43148
rect 4684 43092 4740 43148
rect 35196 43092 35252 43148
rect 35300 43092 35356 43148
rect 35404 43092 35460 43148
rect 19836 42308 19892 42364
rect 19940 42308 19996 42364
rect 20044 42308 20100 42364
rect 50556 42308 50612 42364
rect 50660 42308 50716 42364
rect 50764 42308 50820 42364
rect 4476 41524 4532 41580
rect 4580 41524 4636 41580
rect 4684 41524 4740 41580
rect 35196 41524 35252 41580
rect 35300 41524 35356 41580
rect 35404 41524 35460 41580
rect 19836 40740 19892 40796
rect 19940 40740 19996 40796
rect 20044 40740 20100 40796
rect 50556 40740 50612 40796
rect 50660 40740 50716 40796
rect 50764 40740 50820 40796
rect 40012 40572 40068 40628
rect 40012 40348 40068 40404
rect 4476 39956 4532 40012
rect 4580 39956 4636 40012
rect 4684 39956 4740 40012
rect 35196 39956 35252 40012
rect 35300 39956 35356 40012
rect 35404 39956 35460 40012
rect 5068 39676 5124 39732
rect 19836 39172 19892 39228
rect 19940 39172 19996 39228
rect 20044 39172 20100 39228
rect 50556 39172 50612 39228
rect 50660 39172 50716 39228
rect 50764 39172 50820 39228
rect 9772 38780 9828 38836
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 6076 37996 6132 38052
rect 9772 37660 9828 37716
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 50556 37604 50612 37660
rect 50660 37604 50716 37660
rect 50764 37604 50820 37660
rect 19068 37212 19124 37268
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 6076 36652 6132 36708
rect 19180 36428 19236 36484
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 50556 36036 50612 36092
rect 50660 36036 50716 36092
rect 50764 36036 50820 36092
rect 5068 35868 5124 35924
rect 47068 35532 47124 35588
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 50556 34468 50612 34524
rect 50660 34468 50716 34524
rect 50764 34468 50820 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 50556 32900 50612 32956
rect 50660 32900 50716 32956
rect 50764 32900 50820 32956
rect 6412 32844 6468 32900
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 29932 31948 29988 32004
rect 6412 31388 6468 31444
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 50556 31332 50612 31388
rect 50660 31332 50716 31388
rect 50764 31332 50820 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 47068 30156 47124 30212
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 50556 29764 50612 29820
rect 50660 29764 50716 29820
rect 50764 29764 50820 29820
rect 39676 29484 39732 29540
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19628 28812 19684 28868
rect 47068 28700 47124 28756
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 50556 28196 50612 28252
rect 50660 28196 50716 28252
rect 50764 28196 50820 28252
rect 19628 27692 19684 27748
rect 19516 27468 19572 27524
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 50556 26628 50612 26684
rect 50660 26628 50716 26684
rect 50764 26628 50820 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 32060 25564 32116 25620
rect 37324 25564 37380 25620
rect 19516 25452 19572 25508
rect 31892 25228 31948 25284
rect 37324 25228 37380 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 50556 25060 50612 25116
rect 50660 25060 50716 25116
rect 50764 25060 50820 25116
rect 39676 24556 39732 24612
rect 29932 24332 29988 24388
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 50556 23492 50612 23548
rect 50660 23492 50716 23548
rect 50764 23492 50820 23548
rect 46172 23324 46228 23380
rect 50092 22764 50148 22820
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 5964 22204 6020 22260
rect 41468 22204 41524 22260
rect 49980 21980 50036 22036
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 50556 21924 50612 21980
rect 50660 21924 50716 21980
rect 50764 21924 50820 21980
rect 50092 21868 50148 21924
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 11004 20748 11060 20804
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 50556 20356 50612 20412
rect 50660 20356 50716 20412
rect 50764 20356 50820 20412
rect 39564 20188 39620 20244
rect 43260 20188 43316 20244
rect 25564 19964 25620 20020
rect 39004 19628 39060 19684
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 39788 19516 39844 19572
rect 43260 18844 43316 18900
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 50556 18788 50612 18844
rect 50660 18788 50716 18844
rect 50764 18788 50820 18844
rect 39004 18620 39060 18676
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 50556 17220 50612 17276
rect 50660 17220 50716 17276
rect 50764 17220 50820 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 49980 16156 50036 16212
rect 41468 15708 41524 15764
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 50556 15652 50612 15708
rect 50660 15652 50716 15708
rect 50764 15652 50820 15708
rect 39564 15484 39620 15540
rect 18732 15148 18788 15204
rect 43708 15148 43764 15204
rect 43708 15036 43764 15092
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 50092 14252 50148 14308
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 50556 14084 50612 14140
rect 50660 14084 50716 14140
rect 50764 14084 50820 14140
rect 11004 13916 11060 13972
rect 46172 13916 46228 13972
rect 18732 13580 18788 13636
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 5964 12684 6020 12740
rect 39788 12684 39844 12740
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 50556 12516 50612 12572
rect 50660 12516 50716 12572
rect 50764 12516 50820 12572
rect 25564 12348 25620 12404
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 45388 11228 45444 11284
rect 45612 11228 45668 11284
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 50556 10948 50612 11004
rect 50660 10948 50716 11004
rect 50764 10948 50820 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 50556 9380 50612 9436
rect 50660 9380 50716 9436
rect 50764 9380 50820 9436
rect 45612 8652 45668 8708
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 50556 7812 50612 7868
rect 50660 7812 50716 7868
rect 50764 7812 50820 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 50556 6244 50612 6300
rect 50660 6244 50716 6300
rect 50764 6244 50820 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 50556 4676 50612 4732
rect 50660 4676 50716 4732
rect 50764 4676 50820 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 45388 3388 45444 3444
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
rect 50556 3108 50612 3164
rect 50660 3108 50716 3164
rect 50764 3108 50820 3164
<< metal4 >>
rect 4448 50988 4768 51804
rect 4448 50932 4476 50988
rect 4532 50932 4580 50988
rect 4636 50932 4684 50988
rect 4740 50932 4768 50988
rect 4448 49420 4768 50932
rect 4448 49364 4476 49420
rect 4532 49364 4580 49420
rect 4636 49364 4684 49420
rect 4740 49364 4768 49420
rect 4448 47852 4768 49364
rect 4448 47796 4476 47852
rect 4532 47796 4580 47852
rect 4636 47796 4684 47852
rect 4740 47796 4768 47852
rect 4448 46284 4768 47796
rect 4448 46228 4476 46284
rect 4532 46228 4580 46284
rect 4636 46228 4684 46284
rect 4740 46228 4768 46284
rect 19808 51772 20128 51804
rect 19808 51716 19836 51772
rect 19892 51716 19940 51772
rect 19996 51716 20044 51772
rect 20100 51716 20128 51772
rect 19808 50204 20128 51716
rect 19808 50148 19836 50204
rect 19892 50148 19940 50204
rect 19996 50148 20044 50204
rect 20100 50148 20128 50204
rect 19808 48636 20128 50148
rect 19808 48580 19836 48636
rect 19892 48580 19940 48636
rect 19996 48580 20044 48636
rect 20100 48580 20128 48636
rect 19808 47068 20128 48580
rect 19808 47012 19836 47068
rect 19892 47012 19940 47068
rect 19996 47012 20044 47068
rect 20100 47012 20128 47068
rect 4448 44716 4768 46228
rect 19180 46228 19236 46238
rect 4448 44660 4476 44716
rect 4532 44660 4580 44716
rect 4636 44660 4684 44716
rect 4740 44660 4768 44716
rect 4448 43148 4768 44660
rect 4448 43092 4476 43148
rect 4532 43092 4580 43148
rect 4636 43092 4684 43148
rect 4740 43092 4768 43148
rect 4448 41580 4768 43092
rect 4448 41524 4476 41580
rect 4532 41524 4580 41580
rect 4636 41524 4684 41580
rect 4740 41524 4768 41580
rect 4448 40012 4768 41524
rect 4448 39956 4476 40012
rect 4532 39956 4580 40012
rect 4636 39956 4684 40012
rect 4740 39956 4768 40012
rect 4448 38444 4768 39956
rect 19068 45220 19124 45230
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 5068 39732 5124 39742
rect 5068 35924 5124 39676
rect 9772 38836 9828 38846
rect 6076 38052 6132 38062
rect 6076 36708 6132 37996
rect 9772 37716 9828 38780
rect 9772 37650 9828 37660
rect 19068 37268 19124 45164
rect 19068 37202 19124 37212
rect 6076 36642 6132 36652
rect 19180 36484 19236 46172
rect 19180 36418 19236 36428
rect 19808 45500 20128 47012
rect 19808 45444 19836 45500
rect 19892 45444 19940 45500
rect 19996 45444 20044 45500
rect 20100 45444 20128 45500
rect 19808 43932 20128 45444
rect 19808 43876 19836 43932
rect 19892 43876 19940 43932
rect 19996 43876 20044 43932
rect 20100 43876 20128 43932
rect 19808 42364 20128 43876
rect 19808 42308 19836 42364
rect 19892 42308 19940 42364
rect 19996 42308 20044 42364
rect 20100 42308 20128 42364
rect 19808 40796 20128 42308
rect 19808 40740 19836 40796
rect 19892 40740 19940 40796
rect 19996 40740 20044 40796
rect 20100 40740 20128 40796
rect 19808 39228 20128 40740
rect 19808 39172 19836 39228
rect 19892 39172 19940 39228
rect 19996 39172 20044 39228
rect 20100 39172 20128 39228
rect 19808 37660 20128 39172
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 5068 35858 5124 35868
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 6412 32900 6468 32910
rect 6412 31444 6468 32844
rect 6412 31378 6468 31388
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 35168 50988 35488 51804
rect 35168 50932 35196 50988
rect 35252 50932 35300 50988
rect 35356 50932 35404 50988
rect 35460 50932 35488 50988
rect 35168 49420 35488 50932
rect 35168 49364 35196 49420
rect 35252 49364 35300 49420
rect 35356 49364 35404 49420
rect 35460 49364 35488 49420
rect 35168 47852 35488 49364
rect 35168 47796 35196 47852
rect 35252 47796 35300 47852
rect 35356 47796 35404 47852
rect 35460 47796 35488 47852
rect 35168 46284 35488 47796
rect 50528 51772 50848 51804
rect 50528 51716 50556 51772
rect 50612 51716 50660 51772
rect 50716 51716 50764 51772
rect 50820 51716 50848 51772
rect 50528 50204 50848 51716
rect 50528 50148 50556 50204
rect 50612 50148 50660 50204
rect 50716 50148 50764 50204
rect 50820 50148 50848 50204
rect 50528 48636 50848 50148
rect 50528 48580 50556 48636
rect 50612 48580 50660 48636
rect 50716 48580 50764 48636
rect 50820 48580 50848 48636
rect 50528 47068 50848 48580
rect 50528 47012 50556 47068
rect 50612 47012 50660 47068
rect 50716 47012 50764 47068
rect 50820 47012 50848 47068
rect 35168 46228 35196 46284
rect 35252 46228 35300 46284
rect 35356 46228 35404 46284
rect 35460 46228 35488 46284
rect 35168 44716 35488 46228
rect 35168 44660 35196 44716
rect 35252 44660 35300 44716
rect 35356 44660 35404 44716
rect 35460 44660 35488 44716
rect 35168 43148 35488 44660
rect 35168 43092 35196 43148
rect 35252 43092 35300 43148
rect 35356 43092 35404 43148
rect 35460 43092 35488 43148
rect 35168 41580 35488 43092
rect 35168 41524 35196 41580
rect 35252 41524 35300 41580
rect 35356 41524 35404 41580
rect 35460 41524 35488 41580
rect 35168 40012 35488 41524
rect 47068 46676 47124 46686
rect 40012 40628 40068 40638
rect 40012 40404 40068 40572
rect 40012 40338 40068 40348
rect 35168 39956 35196 40012
rect 35252 39956 35300 40012
rect 35356 39956 35404 40012
rect 35460 39956 35488 40012
rect 35168 38444 35488 39956
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 47068 35588 47124 46620
rect 47068 35522 47124 35532
rect 50528 45500 50848 47012
rect 50528 45444 50556 45500
rect 50612 45444 50660 45500
rect 50716 45444 50764 45500
rect 50820 45444 50848 45500
rect 50528 43932 50848 45444
rect 50528 43876 50556 43932
rect 50612 43876 50660 43932
rect 50716 43876 50764 43932
rect 50820 43876 50848 43932
rect 50528 42364 50848 43876
rect 50528 42308 50556 42364
rect 50612 42308 50660 42364
rect 50716 42308 50764 42364
rect 50820 42308 50848 42364
rect 50528 40796 50848 42308
rect 50528 40740 50556 40796
rect 50612 40740 50660 40796
rect 50716 40740 50764 40796
rect 50820 40740 50848 40796
rect 50528 39228 50848 40740
rect 50528 39172 50556 39228
rect 50612 39172 50660 39228
rect 50716 39172 50764 39228
rect 50820 39172 50848 39228
rect 50528 37660 50848 39172
rect 50528 37604 50556 37660
rect 50612 37604 50660 37660
rect 50716 37604 50764 37660
rect 50820 37604 50848 37660
rect 50528 36092 50848 37604
rect 50528 36036 50556 36092
rect 50612 36036 50660 36092
rect 50716 36036 50764 36092
rect 50820 36036 50848 36092
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19628 28868 19684 28878
rect 19628 27748 19684 28812
rect 19628 27682 19684 27692
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 19516 27524 19572 27534
rect 19516 25508 19572 27468
rect 19516 25442 19572 25452
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 29932 32004 29988 32014
rect 29932 24388 29988 31948
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 50528 34524 50848 36036
rect 50528 34468 50556 34524
rect 50612 34468 50660 34524
rect 50716 34468 50764 34524
rect 50820 34468 50848 34524
rect 50528 32956 50848 34468
rect 50528 32900 50556 32956
rect 50612 32900 50660 32956
rect 50716 32900 50764 32956
rect 50820 32900 50848 32956
rect 50528 31388 50848 32900
rect 50528 31332 50556 31388
rect 50612 31332 50660 31388
rect 50716 31332 50764 31388
rect 50820 31332 50848 31388
rect 47068 30212 47124 30222
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 32060 25620 32116 25630
rect 32060 25498 32116 25564
rect 31948 25442 32116 25498
rect 31948 25318 32004 25442
rect 31892 25284 32004 25318
rect 31948 25262 32004 25284
rect 31892 25218 31948 25228
rect 29932 24322 29988 24332
rect 35168 24332 35488 25844
rect 39676 29540 39732 29550
rect 37324 25620 37380 25630
rect 37324 25284 37380 25564
rect 37324 25218 37380 25228
rect 39676 24612 39732 29484
rect 47068 28756 47124 30156
rect 47068 28690 47124 28700
rect 50528 29820 50848 31332
rect 50528 29764 50556 29820
rect 50612 29764 50660 29820
rect 50716 29764 50764 29820
rect 50820 29764 50848 29820
rect 39676 24546 39732 24556
rect 50528 28252 50848 29764
rect 50528 28196 50556 28252
rect 50612 28196 50660 28252
rect 50716 28196 50764 28252
rect 50820 28196 50848 28252
rect 50528 26684 50848 28196
rect 50528 26628 50556 26684
rect 50612 26628 50660 26684
rect 50716 26628 50764 26684
rect 50820 26628 50848 26684
rect 50528 25116 50848 26628
rect 50528 25060 50556 25116
rect 50612 25060 50660 25116
rect 50716 25060 50764 25116
rect 50820 25060 50848 25116
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 5964 22260 6020 22270
rect 5964 12740 6020 22204
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 11004 20804 11060 20814
rect 11004 13972 11060 20748
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 50528 23548 50848 25060
rect 50528 23492 50556 23548
rect 50612 23492 50660 23548
rect 50716 23492 50764 23548
rect 50820 23492 50848 23548
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 46172 23380 46228 23390
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 11004 13906 11060 13916
rect 18732 15204 18788 15214
rect 18732 13636 18788 15148
rect 18732 13570 18788 13580
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 5964 12674 6020 12684
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 25564 20020 25620 20030
rect 25564 12404 25620 19964
rect 25564 12338 25620 12348
rect 35168 19628 35488 21140
rect 41468 22260 41524 22270
rect 39564 20244 39620 20254
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 39004 19684 39060 19694
rect 39004 18676 39060 19628
rect 39004 18610 39060 18620
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 39564 15540 39620 20188
rect 39564 15474 39620 15484
rect 39788 19572 39844 19582
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 11788 35488 13300
rect 39788 12740 39844 19516
rect 41468 15764 41524 22204
rect 43260 20244 43316 20254
rect 43260 18900 43316 20188
rect 43260 18834 43316 18844
rect 41468 15698 41524 15708
rect 43708 15204 43764 15214
rect 43708 15092 43764 15148
rect 43708 15026 43764 15036
rect 46172 13972 46228 23324
rect 50092 22820 50148 22830
rect 49980 22036 50036 22046
rect 49980 16212 50036 21980
rect 49980 16146 50036 16156
rect 50092 21924 50148 22764
rect 50092 14308 50148 21868
rect 50092 14242 50148 14252
rect 50528 21980 50848 23492
rect 50528 21924 50556 21980
rect 50612 21924 50660 21980
rect 50716 21924 50764 21980
rect 50820 21924 50848 21980
rect 50528 20412 50848 21924
rect 50528 20356 50556 20412
rect 50612 20356 50660 20412
rect 50716 20356 50764 20412
rect 50820 20356 50848 20412
rect 50528 18844 50848 20356
rect 50528 18788 50556 18844
rect 50612 18788 50660 18844
rect 50716 18788 50764 18844
rect 50820 18788 50848 18844
rect 50528 17276 50848 18788
rect 50528 17220 50556 17276
rect 50612 17220 50660 17276
rect 50716 17220 50764 17276
rect 50820 17220 50848 17276
rect 50528 15708 50848 17220
rect 50528 15652 50556 15708
rect 50612 15652 50660 15708
rect 50716 15652 50764 15708
rect 50820 15652 50848 15708
rect 46172 13906 46228 13916
rect 50528 14140 50848 15652
rect 50528 14084 50556 14140
rect 50612 14084 50660 14140
rect 50716 14084 50764 14140
rect 50820 14084 50848 14140
rect 39788 12674 39844 12684
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 50528 12572 50848 14084
rect 50528 12516 50556 12572
rect 50612 12516 50660 12572
rect 50716 12516 50764 12572
rect 50820 12516 50848 12572
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
rect 45388 11284 45444 11294
rect 45388 3444 45444 11228
rect 45612 11284 45668 11294
rect 45612 8708 45668 11228
rect 45612 8642 45668 8652
rect 50528 11004 50848 12516
rect 50528 10948 50556 11004
rect 50612 10948 50660 11004
rect 50716 10948 50764 11004
rect 50820 10948 50848 11004
rect 50528 9436 50848 10948
rect 50528 9380 50556 9436
rect 50612 9380 50660 9436
rect 50716 9380 50764 9436
rect 50820 9380 50848 9436
rect 45388 3378 45444 3388
rect 50528 7868 50848 9380
rect 50528 7812 50556 7868
rect 50612 7812 50660 7868
rect 50716 7812 50764 7868
rect 50820 7812 50848 7868
rect 50528 6300 50848 7812
rect 50528 6244 50556 6300
rect 50612 6244 50660 6300
rect 50716 6244 50764 6300
rect 50820 6244 50848 6300
rect 50528 4732 50848 6244
rect 50528 4676 50556 4732
rect 50612 4676 50660 4732
rect 50716 4676 50764 4732
rect 50820 4676 50848 4732
rect 50528 3164 50848 4676
rect 50528 3108 50556 3164
rect 50612 3108 50660 3164
rect 50716 3108 50764 3164
rect 50820 3108 50848 3164
rect 50528 3076 50848 3108
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0830_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 40096 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0831_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 39088 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0832_
timestamp 1698431365
transform -1 0 49392 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0833_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34496 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0834_
timestamp 1698431365
transform 1 0 34160 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0835_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33824 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0836_
timestamp 1698431365
transform 1 0 33264 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0837_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35056 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai221_4  _0838_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 34832 0 -1 15680
box -86 -86 4902 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0839_
timestamp 1698431365
transform 1 0 40880 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0840_
timestamp 1698431365
transform -1 0 43456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0841_
timestamp 1698431365
transform -1 0 36624 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0842_
timestamp 1698431365
transform -1 0 38640 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0843_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32704 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _0844_
timestamp 1698431365
transform -1 0 36848 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0845_
timestamp 1698431365
transform 1 0 39648 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0846_
timestamp 1698431365
transform -1 0 43008 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0847_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 36960 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_4  _0848_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 42784 0 1 17248
box -86 -86 4566 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0849_
timestamp 1698431365
transform -1 0 40320 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0850_
timestamp 1698431365
transform 1 0 30016 0 1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0851_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38304 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0852_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 38976 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0853_
timestamp 1698431365
transform 1 0 40768 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0854_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44800 0 -1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0855_
timestamp 1698431365
transform 1 0 44912 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _0856_
timestamp 1698431365
transform -1 0 45136 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0857_
timestamp 1698431365
transform -1 0 43792 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0858_
timestamp 1698431365
transform 1 0 43904 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0859_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43680 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _0860_
timestamp 1698431365
transform -1 0 44240 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0861_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 42000 0 -1 20384
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0862_
timestamp 1698431365
transform 1 0 45584 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0863_
timestamp 1698431365
transform -1 0 52976 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0864_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 45472 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0865_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46592 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _0866_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46480 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0867_
timestamp 1698431365
transform 1 0 39760 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0868_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40768 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0869_
timestamp 1698431365
transform 1 0 41440 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0870_
timestamp 1698431365
transform -1 0 44352 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0871_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43680 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0872_
timestamp 1698431365
transform 1 0 46144 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0873_
timestamp 1698431365
transform -1 0 49840 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0874_
timestamp 1698431365
transform 1 0 47488 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0875_
timestamp 1698431365
transform -1 0 49168 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0876_
timestamp 1698431365
transform 1 0 48384 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0877_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0878_
timestamp 1698431365
transform 1 0 47712 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0879_
timestamp 1698431365
transform 1 0 48608 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0880_
timestamp 1698431365
transform 1 0 40768 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0881_
timestamp 1698431365
transform -1 0 41664 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0882_
timestamp 1698431365
transform 1 0 46144 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0883_
timestamp 1698431365
transform -1 0 50400 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0884_
timestamp 1698431365
transform 1 0 48608 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0885_
timestamp 1698431365
transform 1 0 49504 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0886_
timestamp 1698431365
transform 1 0 49280 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0887_
timestamp 1698431365
transform 1 0 50848 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0888_
timestamp 1698431365
transform -1 0 50736 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0889_
timestamp 1698431365
transform 1 0 48608 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0890_
timestamp 1698431365
transform 1 0 49280 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0891_
timestamp 1698431365
transform 1 0 49280 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0892_
timestamp 1698431365
transform 1 0 50736 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0893_
timestamp 1698431365
transform 1 0 47712 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0894_
timestamp 1698431365
transform 1 0 45360 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0895_
timestamp 1698431365
transform 1 0 49056 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0896_
timestamp 1698431365
transform 1 0 49168 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0897_
timestamp 1698431365
transform 1 0 48384 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0898_
timestamp 1698431365
transform -1 0 49952 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0899_
timestamp 1698431365
transform -1 0 50512 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0900_
timestamp 1698431365
transform 1 0 50624 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0901_
timestamp 1698431365
transform 1 0 49616 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0902_
timestamp 1698431365
transform 1 0 46592 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0903_
timestamp 1698431365
transform 1 0 48048 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0904_
timestamp 1698431365
transform 1 0 49168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0905_
timestamp 1698431365
transform -1 0 50624 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0906_
timestamp 1698431365
transform 1 0 50736 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0907_
timestamp 1698431365
transform -1 0 46480 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0908_
timestamp 1698431365
transform 1 0 49392 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0909_
timestamp 1698431365
transform 1 0 48608 0 -1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0910_
timestamp 1698431365
transform -1 0 50400 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0911_
timestamp 1698431365
transform -1 0 50848 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0912_
timestamp 1698431365
transform 1 0 50400 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0913_
timestamp 1698431365
transform -1 0 49168 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0914_
timestamp 1698431365
transform 1 0 47488 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0915_
timestamp 1698431365
transform 1 0 48160 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0916_
timestamp 1698431365
transform -1 0 49280 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0917_
timestamp 1698431365
transform 1 0 48608 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0918_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 53424 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0919_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 46816 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0920_
timestamp 1698431365
transform -1 0 43232 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _0921_
timestamp 1698431365
transform 1 0 44688 0 1 9408
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0922_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46256 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0923_
timestamp 1698431365
transform 1 0 36848 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0924_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 49056 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0925_
timestamp 1698431365
transform 1 0 50624 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0926_
timestamp 1698431365
transform -1 0 53200 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _0927_
timestamp 1698431365
transform -1 0 50064 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0928_
timestamp 1698431365
transform -1 0 49952 0 -1 9408
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0929_
timestamp 1698431365
transform -1 0 45920 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0930_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48496 0 1 7840
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0931_
timestamp 1698431365
transform 1 0 50400 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0932_
timestamp 1698431365
transform -1 0 48832 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _0933_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 49728 0 -1 7840
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0934_
timestamp 1698431365
transform -1 0 48384 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0935_
timestamp 1698431365
transform 1 0 47936 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _0936_
timestamp 1698431365
transform 1 0 49280 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0937_
timestamp 1698431365
transform 1 0 49728 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0938_
timestamp 1698431365
transform -1 0 45696 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _0939_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44688 0 1 7840
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _0940_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44240 0 -1 7840
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0941_
timestamp 1698431365
transform 1 0 44688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _0942_
timestamp 1698431365
transform 1 0 40096 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _0943_
timestamp 1698431365
transform -1 0 41664 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0944_
timestamp 1698431365
transform 1 0 41888 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0945_
timestamp 1698431365
transform -1 0 42112 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _0946_
timestamp 1698431365
transform 1 0 45696 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0947_
timestamp 1698431365
transform 1 0 41664 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _0948_
timestamp 1698431365
transform 1 0 41664 0 1 6272
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0949_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41664 0 -1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0950_
timestamp 1698431365
transform 1 0 44128 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0951_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43008 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0952_
timestamp 1698431365
transform 1 0 24192 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0953_
timestamp 1698431365
transform 1 0 25312 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0954_
timestamp 1698431365
transform 1 0 25536 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0955_
timestamp 1698431365
transform -1 0 27776 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0956_
timestamp 1698431365
transform -1 0 36512 0 -1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0957_
timestamp 1698431365
transform 1 0 32928 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0958_
timestamp 1698431365
transform -1 0 44240 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0959_
timestamp 1698431365
transform -1 0 43008 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _0960_
timestamp 1698431365
transform -1 0 40544 0 -1 9408
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0961_
timestamp 1698431365
transform 1 0 39536 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0962_
timestamp 1698431365
transform 1 0 41776 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _0963_
timestamp 1698431365
transform -1 0 41440 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0964_
timestamp 1698431365
transform -1 0 42784 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0965_
timestamp 1698431365
transform -1 0 43568 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0966_
timestamp 1698431365
transform 1 0 45920 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0967_
timestamp 1698431365
transform -1 0 42448 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0968_
timestamp 1698431365
transform -1 0 43120 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0969_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41888 0 -1 15680
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _0970_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 41104 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0971_
timestamp 1698431365
transform 1 0 43344 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0972_
timestamp 1698431365
transform 1 0 44240 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0973_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 41664 0 -1 15680
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0974_
timestamp 1698431365
transform 1 0 40432 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _0975_
timestamp 1698431365
transform -1 0 42560 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0976_
timestamp 1698431365
transform -1 0 38528 0 1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0977_
timestamp 1698431365
transform 1 0 37968 0 1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0978_
timestamp 1698431365
transform -1 0 38976 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0979_
timestamp 1698431365
transform -1 0 38640 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _0980_
timestamp 1698431365
transform -1 0 38976 0 1 15680
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _0981_
timestamp 1698431365
transform 1 0 35056 0 -1 14112
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0982_
timestamp 1698431365
transform -1 0 36512 0 1 12544
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0983_
timestamp 1698431365
transform 1 0 36176 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0984_
timestamp 1698431365
transform 1 0 30464 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _0985_
timestamp 1698431365
transform -1 0 36064 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0986_
timestamp 1698431365
transform -1 0 33376 0 1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _0987_
timestamp 1698431365
transform -1 0 32816 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _0988_
timestamp 1698431365
transform -1 0 32032 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0989_
timestamp 1698431365
transform -1 0 31696 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _0990_
timestamp 1698431365
transform 1 0 31696 0 -1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _0991_
timestamp 1698431365
transform 1 0 33488 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _0992_
timestamp 1698431365
transform -1 0 36400 0 1 9408
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0993_
timestamp 1698431365
transform -1 0 32704 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _0994_
timestamp 1698431365
transform 1 0 25760 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0995_
timestamp 1698431365
transform -1 0 32144 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _0996_
timestamp 1698431365
transform -1 0 34048 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _0997_
timestamp 1698431365
transform 1 0 35280 0 -1 9408
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _0998_
timestamp 1698431365
transform -1 0 33488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _0999_
timestamp 1698431365
transform 1 0 39760 0 1 9408
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1000_
timestamp 1698431365
transform -1 0 30688 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1001_
timestamp 1698431365
transform 1 0 29792 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1002_
timestamp 1698431365
transform -1 0 38528 0 1 6272
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1003_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 48384 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1004_
timestamp 1698431365
transform -1 0 38528 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1005_
timestamp 1698431365
transform -1 0 31808 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1006_
timestamp 1698431365
transform 1 0 35952 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1007_
timestamp 1698431365
transform 1 0 31584 0 1 6272
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1008_
timestamp 1698431365
transform 1 0 27328 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1009_
timestamp 1698431365
transform -1 0 26320 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1010_
timestamp 1698431365
transform -1 0 25648 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1011_
timestamp 1698431365
transform 1 0 27104 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1012_
timestamp 1698431365
transform 1 0 27328 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1013_
timestamp 1698431365
transform -1 0 27104 0 1 6272
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1014_
timestamp 1698431365
transform 1 0 27440 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1015_
timestamp 1698431365
transform -1 0 27440 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1016_
timestamp 1698431365
transform -1 0 25760 0 -1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1017_
timestamp 1698431365
transform 1 0 21168 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1018_
timestamp 1698431365
transform -1 0 24528 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1019_
timestamp 1698431365
transform 1 0 21392 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1020_
timestamp 1698431365
transform -1 0 22400 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1021_
timestamp 1698431365
transform -1 0 22512 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1022_
timestamp 1698431365
transform -1 0 21280 0 -1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1023_
timestamp 1698431365
transform -1 0 24416 0 -1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1024_
timestamp 1698431365
transform -1 0 22400 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1025_
timestamp 1698431365
transform -1 0 22288 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1026_
timestamp 1698431365
transform -1 0 23072 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1027_
timestamp 1698431365
transform 1 0 21168 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1028_
timestamp 1698431365
transform 1 0 22624 0 1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1029_
timestamp 1698431365
transform -1 0 23856 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1030_
timestamp 1698431365
transform -1 0 23632 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1031_
timestamp 1698431365
transform -1 0 25872 0 -1 9408
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1032_
timestamp 1698431365
transform -1 0 25648 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1033_
timestamp 1698431365
transform 1 0 22512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1034_
timestamp 1698431365
transform 1 0 25088 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1035_
timestamp 1698431365
transform 1 0 38528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _1036_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37744 0 1 4704
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1037_
timestamp 1698431365
transform 1 0 36960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1038_
timestamp 1698431365
transform 1 0 25760 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1039_
timestamp 1698431365
transform -1 0 44128 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1040_
timestamp 1698431365
transform -1 0 44016 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1041_
timestamp 1698431365
transform -1 0 41440 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1042_
timestamp 1698431365
transform -1 0 36064 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1043_
timestamp 1698431365
transform -1 0 33936 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1044_
timestamp 1698431365
transform -1 0 34944 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1045_
timestamp 1698431365
transform 1 0 34832 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1046_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 33936 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1047_
timestamp 1698431365
transform -1 0 34160 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1048_
timestamp 1698431365
transform 1 0 25424 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1049_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 43344 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1050_
timestamp 1698431365
transform -1 0 31920 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1051_
timestamp 1698431365
transform 1 0 32144 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1052_
timestamp 1698431365
transform -1 0 34048 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1053_
timestamp 1698431365
transform -1 0 33488 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1054_
timestamp 1698431365
transform -1 0 47488 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1055_
timestamp 1698431365
transform -1 0 30688 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1056_
timestamp 1698431365
transform -1 0 29904 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1057_
timestamp 1698431365
transform 1 0 29904 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1058_
timestamp 1698431365
transform -1 0 46704 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1059_
timestamp 1698431365
transform 1 0 30688 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1060_
timestamp 1698431365
transform 1 0 30128 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1061_
timestamp 1698431365
transform 1 0 30688 0 1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1062_
timestamp 1698431365
transform -1 0 46592 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1063_
timestamp 1698431365
transform -1 0 31472 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1064_
timestamp 1698431365
transform -1 0 34832 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1065_
timestamp 1698431365
transform 1 0 29568 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1066_
timestamp 1698431365
transform 1 0 30128 0 1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1067_
timestamp 1698431365
transform -1 0 34496 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1068_
timestamp 1698431365
transform -1 0 46928 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1069_
timestamp 1698431365
transform -1 0 30128 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1070_
timestamp 1698431365
transform -1 0 30688 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1071_
timestamp 1698431365
transform -1 0 30128 0 1 28224
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1072_
timestamp 1698431365
transform -1 0 47824 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1073_
timestamp 1698431365
transform -1 0 30016 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1074_
timestamp 1698431365
transform -1 0 29568 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1075_
timestamp 1698431365
transform 1 0 29232 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1076_
timestamp 1698431365
transform -1 0 46928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1077_
timestamp 1698431365
transform -1 0 31360 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1078_
timestamp 1698431365
transform -1 0 31136 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1079_
timestamp 1698431365
transform -1 0 30912 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1080_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 46704 0 1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1081_
timestamp 1698431365
transform 1 0 47712 0 -1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1082_
timestamp 1698431365
transform -1 0 41440 0 1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1083_
timestamp 1698431365
transform 1 0 49280 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1084_
timestamp 1698431365
transform 1 0 44688 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1085_
timestamp 1698431365
transform 1 0 47712 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1086_
timestamp 1698431365
transform -1 0 37744 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1087_
timestamp 1698431365
transform 1 0 41328 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1088_
timestamp 1698431365
transform 1 0 43568 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1089_
timestamp 1698431365
transform -1 0 42672 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1090_
timestamp 1698431365
transform -1 0 39312 0 -1 34496
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1091_
timestamp 1698431365
transform 1 0 41440 0 1 26656
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _1092_
timestamp 1698431365
transform -1 0 44912 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1093_
timestamp 1698431365
transform -1 0 25872 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1094_
timestamp 1698431365
transform 1 0 37408 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1095_
timestamp 1698431365
transform 1 0 38976 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1096_
timestamp 1698431365
transform -1 0 44576 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1097_
timestamp 1698431365
transform 1 0 41888 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1098_
timestamp 1698431365
transform 1 0 42336 0 -1 23520
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1099_
timestamp 1698431365
transform 1 0 25648 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1100_
timestamp 1698431365
transform -1 0 43120 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1101_
timestamp 1698431365
transform -1 0 42000 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1102_
timestamp 1698431365
transform 1 0 42224 0 1 25088
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1103_
timestamp 1698431365
transform -1 0 37744 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1104_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 37520 0 -1 23520
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1105_
timestamp 1698431365
transform 1 0 44576 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _1106_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1107_
timestamp 1698431365
transform 1 0 50064 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1108_
timestamp 1698431365
transform -1 0 43568 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1109_
timestamp 1698431365
transform -1 0 39648 0 1 34496
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1110_
timestamp 1698431365
transform -1 0 38752 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1111_
timestamp 1698431365
transform -1 0 44240 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1112_
timestamp 1698431365
transform 1 0 37520 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1113_
timestamp 1698431365
transform 1 0 38640 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1114_
timestamp 1698431365
transform 1 0 37968 0 -1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1115_
timestamp 1698431365
transform -1 0 49504 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1116_
timestamp 1698431365
transform 1 0 45248 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi222_2  _1117_
timestamp 1698431365
transform 1 0 36400 0 -1 36064
box -86 -86 2886 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1118_
timestamp 1698431365
transform 1 0 28672 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1119_
timestamp 1698431365
transform 1 0 38640 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_2  _1120_
timestamp 1698431365
transform -1 0 41328 0 1 25088
box -86 -86 2662 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1121_
timestamp 1698431365
transform 1 0 42000 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1122_
timestamp 1698431365
transform -1 0 49504 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1123_
timestamp 1698431365
transform 1 0 45920 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1124_
timestamp 1698431365
transform 1 0 48608 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1125_
timestamp 1698431365
transform 1 0 44688 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1126_
timestamp 1698431365
transform -1 0 24864 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1127_
timestamp 1698431365
transform 1 0 23856 0 1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1128_
timestamp 1698431365
transform 1 0 36064 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1129_
timestamp 1698431365
transform 1 0 42896 0 -1 31360
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1130_
timestamp 1698431365
transform -1 0 50848 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1131_
timestamp 1698431365
transform 1 0 50848 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1132_
timestamp 1698431365
transform -1 0 44128 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1133_
timestamp 1698431365
transform -1 0 25088 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1134_
timestamp 1698431365
transform 1 0 23184 0 1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1135_
timestamp 1698431365
transform -1 0 36400 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1136_
timestamp 1698431365
transform -1 0 36960 0 -1 28224
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1137_
timestamp 1698431365
transform 1 0 42784 0 -1 32928
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1138_
timestamp 1698431365
transform -1 0 50736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1139_
timestamp 1698431365
transform -1 0 50176 0 -1 34496
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1140_
timestamp 1698431365
transform 1 0 43568 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1141_
timestamp 1698431365
transform -1 0 24528 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1142_
timestamp 1698431365
transform -1 0 35952 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1143_
timestamp 1698431365
transform 1 0 42448 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1144_
timestamp 1698431365
transform -1 0 50960 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1145_
timestamp 1698431365
transform 1 0 50960 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1146_
timestamp 1698431365
transform 1 0 48608 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1147_
timestamp 1698431365
transform -1 0 42896 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1148_
timestamp 1698431365
transform 1 0 23184 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1149_
timestamp 1698431365
transform -1 0 36288 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1150_
timestamp 1698431365
transform 1 0 41552 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1151_
timestamp 1698431365
transform -1 0 49392 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1152_
timestamp 1698431365
transform 1 0 49504 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1153_
timestamp 1698431365
transform -1 0 40096 0 -1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_2  _1154_
timestamp 1698431365
transform 1 0 24864 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1155_
timestamp 1698431365
transform -1 0 36624 0 -1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1156_
timestamp 1698431365
transform 1 0 38640 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1157_
timestamp 1698431365
transform -1 0 51184 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1158_
timestamp 1698431365
transform 1 0 51184 0 1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1159_
timestamp 1698431365
transform 1 0 32704 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1160_
timestamp 1698431365
transform 1 0 14784 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1161_
timestamp 1698431365
transform -1 0 19936 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1162_
timestamp 1698431365
transform 1 0 17248 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1163_
timestamp 1698431365
transform -1 0 19712 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1164_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 18928 0 1 37632
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1165_
timestamp 1698431365
transform 1 0 16576 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1166_
timestamp 1698431365
transform -1 0 21392 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1167_
timestamp 1698431365
transform 1 0 18256 0 1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1168_
timestamp 1698431365
transform 1 0 15680 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1169_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 18928 0 1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1170_
timestamp 1698431365
transform -1 0 20048 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1171_
timestamp 1698431365
transform 1 0 31248 0 -1 40768
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1172_
timestamp 1698431365
transform -1 0 34496 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1173_
timestamp 1698431365
transform 1 0 29344 0 -1 39200
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1174_
timestamp 1698431365
transform 1 0 30240 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1175_
timestamp 1698431365
transform 1 0 30688 0 -1 39200
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1176_
timestamp 1698431365
transform 1 0 27440 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1177_
timestamp 1698431365
transform 1 0 25088 0 -1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1178_
timestamp 1698431365
transform 1 0 27440 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1179_
timestamp 1698431365
transform 1 0 25312 0 1 37632
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1180_
timestamp 1698431365
transform 1 0 27776 0 -1 37632
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1181_
timestamp 1698431365
transform 1 0 31808 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1182_
timestamp 1698431365
transform 1 0 32928 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1183_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 48608 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1184_
timestamp 1698431365
transform 1 0 33264 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _1185_
timestamp 1698431365
transform -1 0 37632 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1186_
timestamp 1698431365
transform 1 0 38640 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1187_
timestamp 1698431365
transform 1 0 46592 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1188_
timestamp 1698431365
transform -1 0 47264 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1189_
timestamp 1698431365
transform 1 0 48608 0 1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1190_
timestamp 1698431365
transform 1 0 49168 0 1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1191_
timestamp 1698431365
transform 1 0 50624 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1192_
timestamp 1698431365
transform 1 0 49728 0 -1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1193_
timestamp 1698431365
transform 1 0 48608 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1194_
timestamp 1698431365
transform -1 0 50848 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1195_
timestamp 1698431365
transform 1 0 51072 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1196_
timestamp 1698431365
transform 1 0 48944 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1197_
timestamp 1698431365
transform -1 0 50288 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1198_
timestamp 1698431365
transform -1 0 49392 0 1 48608
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1199_
timestamp 1698431365
transform -1 0 48384 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1200_
timestamp 1698431365
transform 1 0 48272 0 1 43904
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1201_
timestamp 1698431365
transform 1 0 48944 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1202_
timestamp 1698431365
transform 1 0 50400 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1203_
timestamp 1698431365
transform 1 0 25984 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1204_
timestamp 1698431365
transform 1 0 37408 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1205_
timestamp 1698431365
transform 1 0 39200 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1206_
timestamp 1698431365
transform 1 0 38080 0 -1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1207_
timestamp 1698431365
transform -1 0 25984 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1208_
timestamp 1698431365
transform 1 0 23184 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1209_
timestamp 1698431365
transform 1 0 25312 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1210_
timestamp 1698431365
transform -1 0 20160 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1211_
timestamp 1698431365
transform -1 0 19936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1212_
timestamp 1698431365
transform -1 0 26208 0 -1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1213_
timestamp 1698431365
transform 1 0 25424 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1214_
timestamp 1698431365
transform -1 0 25536 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1215_
timestamp 1698431365
transform -1 0 22736 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1216_
timestamp 1698431365
transform 1 0 24416 0 1 34496
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1217_
timestamp 1698431365
transform 1 0 25424 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1218_
timestamp 1698431365
transform -1 0 23744 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1219_
timestamp 1698431365
transform 1 0 22064 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1220_
timestamp 1698431365
transform 1 0 22624 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1221_
timestamp 1698431365
transform -1 0 23296 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1222_
timestamp 1698431365
transform 1 0 20384 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1223_
timestamp 1698431365
transform -1 0 21952 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1224_
timestamp 1698431365
transform 1 0 21168 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1225_
timestamp 1698431365
transform -1 0 23408 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1226_
timestamp 1698431365
transform 1 0 20160 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1227_
timestamp 1698431365
transform 1 0 20384 0 1 29792
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1228_
timestamp 1698431365
transform 1 0 21168 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1229_
timestamp 1698431365
transform -1 0 19600 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1230_
timestamp 1698431365
transform 1 0 19376 0 1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1231_
timestamp 1698431365
transform 1 0 19600 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1232_
timestamp 1698431365
transform -1 0 20832 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1233_
timestamp 1698431365
transform -1 0 20048 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1234_
timestamp 1698431365
transform 1 0 19376 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1235_
timestamp 1698431365
transform -1 0 23184 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1236_
timestamp 1698431365
transform 1 0 22064 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1237_
timestamp 1698431365
transform 1 0 23408 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1238_
timestamp 1698431365
transform 1 0 22288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1239_
timestamp 1698431365
transform -1 0 32480 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1240_
timestamp 1698431365
transform -1 0 31472 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1241_
timestamp 1698431365
transform -1 0 31360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1242_
timestamp 1698431365
transform 1 0 36848 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1243_
timestamp 1698431365
transform 1 0 34944 0 1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1244_
timestamp 1698431365
transform 1 0 31024 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1245_
timestamp 1698431365
transform 1 0 31696 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1246_
timestamp 1698431365
transform 1 0 33040 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1247_
timestamp 1698431365
transform -1 0 35168 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1248_
timestamp 1698431365
transform -1 0 34608 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1249_
timestamp 1698431365
transform 1 0 34160 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1250_
timestamp 1698431365
transform 1 0 34720 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1251_
timestamp 1698431365
transform -1 0 32032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1252_
timestamp 1698431365
transform 1 0 31360 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1253_
timestamp 1698431365
transform 1 0 32368 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1254_
timestamp 1698431365
transform 1 0 27888 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1255_
timestamp 1698431365
transform -1 0 30800 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1256_
timestamp 1698431365
transform -1 0 28672 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1257_
timestamp 1698431365
transform -1 0 28224 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1258_
timestamp 1698431365
transform -1 0 29680 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1259_
timestamp 1698431365
transform -1 0 28448 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1260_
timestamp 1698431365
transform 1 0 33824 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1261_
timestamp 1698431365
transform 1 0 33152 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1262_
timestamp 1698431365
transform -1 0 29008 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1263_
timestamp 1698431365
transform -1 0 29568 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1264_
timestamp 1698431365
transform -1 0 27776 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1265_
timestamp 1698431365
transform -1 0 27552 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1266_
timestamp 1698431365
transform -1 0 32480 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1267_
timestamp 1698431365
transform 1 0 28112 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1268_
timestamp 1698431365
transform 1 0 33936 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1269_
timestamp 1698431365
transform 1 0 33264 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1270_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 35504 0 -1 45472
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1271_
timestamp 1698431365
transform 1 0 23856 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1272_
timestamp 1698431365
transform 1 0 26768 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1273_
timestamp 1698431365
transform -1 0 27552 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1274_
timestamp 1698431365
transform 1 0 29568 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1275_
timestamp 1698431365
transform 1 0 21952 0 1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1276_
timestamp 1698431365
transform 1 0 25872 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1277_
timestamp 1698431365
transform 1 0 25872 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1278_
timestamp 1698431365
transform 1 0 33824 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1279_
timestamp 1698431365
transform -1 0 33824 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1280_
timestamp 1698431365
transform -1 0 23744 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1281_
timestamp 1698431365
transform 1 0 25536 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1282_
timestamp 1698431365
transform -1 0 21392 0 -1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1283_
timestamp 1698431365
transform 1 0 20944 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1284_
timestamp 1698431365
transform -1 0 25872 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1285_
timestamp 1698431365
transform -1 0 28672 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1286_
timestamp 1698431365
transform 1 0 15904 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1287_
timestamp 1698431365
transform -1 0 24192 0 1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1288_
timestamp 1698431365
transform -1 0 23072 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1289_
timestamp 1698431365
transform 1 0 23184 0 -1 42336
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1290_
timestamp 1698431365
transform -1 0 26880 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1291_
timestamp 1698431365
transform 1 0 26208 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1292_
timestamp 1698431365
transform -1 0 24640 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1293_
timestamp 1698431365
transform 1 0 24080 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1294_
timestamp 1698431365
transform -1 0 23744 0 1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1295_
timestamp 1698431365
transform 1 0 22624 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1296_
timestamp 1698431365
transform 1 0 22400 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1297_
timestamp 1698431365
transform -1 0 22400 0 1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1298_
timestamp 1698431365
transform 1 0 19936 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1299_
timestamp 1698431365
transform 1 0 22848 0 -1 40768
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _1300_
timestamp 1698431365
transform -1 0 24976 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1301_
timestamp 1698431365
transform 1 0 23632 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1302_
timestamp 1698431365
transform -1 0 38640 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1303_
timestamp 1698431365
transform -1 0 25984 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1304_
timestamp 1698431365
transform -1 0 25312 0 1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1305_
timestamp 1698431365
transform 1 0 24528 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1306_
timestamp 1698431365
transform 1 0 23072 0 -1 50176
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1307_
timestamp 1698431365
transform 1 0 23856 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1308_
timestamp 1698431365
transform -1 0 40320 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1309_
timestamp 1698431365
transform -1 0 31584 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1310_
timestamp 1698431365
transform 1 0 23856 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1311_
timestamp 1698431365
transform 1 0 25088 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1312_
timestamp 1698431365
transform 1 0 31584 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1313_
timestamp 1698431365
transform -1 0 27552 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1314_
timestamp 1698431365
transform -1 0 27328 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1315_
timestamp 1698431365
transform 1 0 27216 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1316_
timestamp 1698431365
transform -1 0 25648 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1317_
timestamp 1698431365
transform 1 0 25648 0 1 47040
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1318_
timestamp 1698431365
transform -1 0 28448 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1319_
timestamp 1698431365
transform 1 0 27104 0 -1 50176
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1320_
timestamp 1698431365
transform -1 0 27440 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1321_
timestamp 1698431365
transform 1 0 26320 0 -1 50176
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1322_
timestamp 1698431365
transform 1 0 27104 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1323_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 29904 0 -1 47040
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1324_
timestamp 1698431365
transform 1 0 21616 0 1 45472
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1325_
timestamp 1698431365
transform -1 0 34048 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1326_
timestamp 1698431365
transform 1 0 19376 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1327_
timestamp 1698431365
transform 1 0 20272 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1328_
timestamp 1698431365
transform 1 0 21952 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1329_
timestamp 1698431365
transform -1 0 21952 0 -1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1330_
timestamp 1698431365
transform 1 0 31472 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1331_
timestamp 1698431365
transform -1 0 19040 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1332_
timestamp 1698431365
transform -1 0 18704 0 1 48608
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1333_
timestamp 1698431365
transform -1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1334_
timestamp 1698431365
transform -1 0 20048 0 1 48608
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1335_
timestamp 1698431365
transform 1 0 10752 0 -1 43904
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1336_
timestamp 1698431365
transform -1 0 18144 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1337_
timestamp 1698431365
transform -1 0 19824 0 1 47040
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1338_
timestamp 1698431365
transform 1 0 17920 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1339_
timestamp 1698431365
transform 1 0 18816 0 -1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1340_
timestamp 1698431365
transform -1 0 18928 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1341_
timestamp 1698431365
transform -1 0 18032 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1342_
timestamp 1698431365
transform 1 0 19264 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1343_
timestamp 1698431365
transform 1 0 19712 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1344_
timestamp 1698431365
transform 1 0 19936 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1345_
timestamp 1698431365
transform 1 0 18256 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1346_
timestamp 1698431365
transform 1 0 18704 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1347_
timestamp 1698431365
transform 1 0 20720 0 -1 47040
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1348_
timestamp 1698431365
transform 1 0 11984 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _1349_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 15344 0 1 45472
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1350_
timestamp 1698431365
transform -1 0 12544 0 -1 47040
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1351_
timestamp 1698431365
transform 1 0 11872 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1352_
timestamp 1698431365
transform -1 0 11984 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1353_
timestamp 1698431365
transform 1 0 12992 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1354_
timestamp 1698431365
transform -1 0 15344 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _1355_
timestamp 1698431365
transform 1 0 13888 0 -1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1356_
timestamp 1698431365
transform -1 0 14672 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1357_
timestamp 1698431365
transform 1 0 12208 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1358_
timestamp 1698431365
transform 1 0 13888 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _1359_
timestamp 1698431365
transform 1 0 13664 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1360_
timestamp 1698431365
transform -1 0 15344 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1361_
timestamp 1698431365
transform -1 0 14784 0 -1 43904
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1362_
timestamp 1698431365
transform -1 0 12880 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1363_
timestamp 1698431365
transform -1 0 12320 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1364_
timestamp 1698431365
transform -1 0 15680 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1365_
timestamp 1698431365
transform -1 0 14784 0 -1 42336
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1366_
timestamp 1698431365
transform 1 0 14560 0 1 42336
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1367_
timestamp 1698431365
transform 1 0 14224 0 1 40768
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1368_
timestamp 1698431365
transform -1 0 49728 0 -1 45472
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1369_
timestamp 1698431365
transform 1 0 35504 0 -1 45472
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1370_
timestamp 1698431365
transform 1 0 37744 0 1 45472
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1371_
timestamp 1698431365
transform -1 0 40544 0 -1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1372_
timestamp 1698431365
transform -1 0 36624 0 1 43904
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1373_
timestamp 1698431365
transform -1 0 40096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1374_
timestamp 1698431365
transform 1 0 37856 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1375_
timestamp 1698431365
transform 1 0 38192 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1376_
timestamp 1698431365
transform -1 0 38192 0 -1 50176
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1377_
timestamp 1698431365
transform -1 0 35616 0 1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1378_
timestamp 1698431365
transform -1 0 42672 0 -1 48608
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1379_
timestamp 1698431365
transform -1 0 41776 0 1 48608
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1380_
timestamp 1698431365
transform 1 0 41664 0 -1 50176
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1381_
timestamp 1698431365
transform 1 0 40096 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1382_
timestamp 1698431365
transform -1 0 42448 0 1 47040
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1383_
timestamp 1698431365
transform 1 0 42560 0 1 47040
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1384_
timestamp 1698431365
transform -1 0 43680 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1385_
timestamp 1698431365
transform 1 0 43680 0 1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1386_
timestamp 1698431365
transform 1 0 41664 0 1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1387_
timestamp 1698431365
transform 1 0 42784 0 -1 45472
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_2  _1388_
timestamp 1698431365
transform -1 0 25760 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1389_
timestamp 1698431365
transform 1 0 40768 0 -1 45472
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1390_
timestamp 1698431365
transform -1 0 41440 0 -1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1391_
timestamp 1698431365
transform 1 0 38528 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1392_
timestamp 1698431365
transform 1 0 36848 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1393_
timestamp 1698431365
transform 1 0 32928 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1394_
timestamp 1698431365
transform 1 0 38304 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1395_
timestamp 1698431365
transform -1 0 39872 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1396_
timestamp 1698431365
transform -1 0 29680 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1397_
timestamp 1698431365
transform 1 0 14224 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1398_
timestamp 1698431365
transform 1 0 15680 0 -1 25088
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _1399_
timestamp 1698431365
transform 1 0 17696 0 -1 25088
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1400_
timestamp 1698431365
transform -1 0 17024 0 -1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1401_
timestamp 1698431365
transform 1 0 15120 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _1402_
timestamp 1698431365
transform 1 0 16016 0 1 29792
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1403_
timestamp 1698431365
transform 1 0 17248 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1404_
timestamp 1698431365
transform 1 0 15680 0 -1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1405_
timestamp 1698431365
transform 1 0 16240 0 1 28224
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1406_
timestamp 1698431365
transform 1 0 14336 0 -1 29792
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_4  _1407_
timestamp 1698431365
transform 1 0 17248 0 -1 28224
box -86 -86 4230 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _1408_
timestamp 1698431365
transform 1 0 15904 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1409_
timestamp 1698431365
transform -1 0 9184 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1410_
timestamp 1698431365
transform 1 0 17808 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1411_
timestamp 1698431365
transform 1 0 18368 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1412_
timestamp 1698431365
transform 1 0 17360 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1413_
timestamp 1698431365
transform 1 0 17472 0 -1 31360
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _1414_
timestamp 1698431365
transform 1 0 18704 0 -1 32928
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1415_
timestamp 1698431365
transform 1 0 14112 0 1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1416_
timestamp 1698431365
transform 1 0 14448 0 1 36064
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1417_
timestamp 1698431365
transform 1 0 13888 0 1 34496
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1418_
timestamp 1698431365
transform 1 0 13216 0 -1 32928
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _1419_
timestamp 1698431365
transform 1 0 14672 0 -1 32928
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1420_
timestamp 1698431365
transform 1 0 15904 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1421_
timestamp 1698431365
transform -1 0 8176 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1422_
timestamp 1698431365
transform 1 0 4480 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1423_
timestamp 1698431365
transform -1 0 41440 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _1424_
timestamp 1698431365
transform -1 0 40432 0 -1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1425_
timestamp 1698431365
transform -1 0 9072 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1426_
timestamp 1698431365
transform 1 0 7168 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1427_
timestamp 1698431365
transform 1 0 4368 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1428_
timestamp 1698431365
transform 1 0 4704 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1429_
timestamp 1698431365
transform 1 0 5488 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1430_
timestamp 1698431365
transform -1 0 10640 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1431_
timestamp 1698431365
transform 1 0 14336 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1432_
timestamp 1698431365
transform -1 0 14336 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1433_
timestamp 1698431365
transform 1 0 7840 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1434_
timestamp 1698431365
transform -1 0 7392 0 -1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1435_
timestamp 1698431365
transform -1 0 8512 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1436_
timestamp 1698431365
transform -1 0 2800 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1437_
timestamp 1698431365
transform 1 0 4816 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1438_
timestamp 1698431365
transform -1 0 40544 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1439_
timestamp 1698431365
transform -1 0 15680 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1440_
timestamp 1698431365
transform -1 0 10752 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1441_
timestamp 1698431365
transform 1 0 5824 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1442_
timestamp 1698431365
transform 1 0 6832 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1443_
timestamp 1698431365
transform -1 0 7392 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1444_
timestamp 1698431365
transform 1 0 7504 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1445_
timestamp 1698431365
transform -1 0 30912 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1446_
timestamp 1698431365
transform -1 0 7056 0 -1 14112
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _1447_
timestamp 1698431365
transform 1 0 4816 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1448_
timestamp 1698431365
transform 1 0 6160 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1449_
timestamp 1698431365
transform -1 0 10080 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _1450_
timestamp 1698431365
transform -1 0 6944 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1451_
timestamp 1698431365
transform 1 0 6384 0 1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1452_
timestamp 1698431365
transform 1 0 4816 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1453_
timestamp 1698431365
transform 1 0 5488 0 1 12544
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1454_
timestamp 1698431365
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1455_
timestamp 1698431365
transform -1 0 12656 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1456_
timestamp 1698431365
transform -1 0 11536 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1457_
timestamp 1698431365
transform -1 0 6720 0 1 10976
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1458_
timestamp 1698431365
transform -1 0 9520 0 1 10976
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1459_
timestamp 1698431365
transform 1 0 7056 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1460_
timestamp 1698431365
transform -1 0 12208 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1461_
timestamp 1698431365
transform 1 0 7728 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1462_
timestamp 1698431365
transform -1 0 8512 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1463_
timestamp 1698431365
transform -1 0 8960 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1464_
timestamp 1698431365
transform 1 0 12992 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1465_
timestamp 1698431365
transform 1 0 10864 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1466_
timestamp 1698431365
transform 1 0 10528 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1467_
timestamp 1698431365
transform 1 0 9744 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1468_
timestamp 1698431365
transform -1 0 11872 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1469_
timestamp 1698431365
transform -1 0 14224 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1470_
timestamp 1698431365
transform -1 0 16352 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1471_
timestamp 1698431365
transform -1 0 15008 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1472_
timestamp 1698431365
transform 1 0 11984 0 -1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1473_
timestamp 1698431365
transform -1 0 12992 0 -1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1474_
timestamp 1698431365
transform -1 0 16240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1475_
timestamp 1698431365
transform 1 0 12656 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1476_
timestamp 1698431365
transform -1 0 14336 0 -1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1477_
timestamp 1698431365
transform 1 0 13776 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1478_
timestamp 1698431365
transform -1 0 19040 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1479_
timestamp 1698431365
transform 1 0 13888 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1480_
timestamp 1698431365
transform -1 0 19488 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1481_
timestamp 1698431365
transform 1 0 17136 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1482_
timestamp 1698431365
transform 1 0 15344 0 1 12544
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1483_
timestamp 1698431365
transform -1 0 16576 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1484_
timestamp 1698431365
transform 1 0 15008 0 1 10976
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1485_
timestamp 1698431365
transform -1 0 20944 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1486_
timestamp 1698431365
transform 1 0 12096 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1487_
timestamp 1698431365
transform 1 0 16464 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1488_
timestamp 1698431365
transform 1 0 19264 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1489_
timestamp 1698431365
transform 1 0 18144 0 -1 14112
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1490_
timestamp 1698431365
transform 1 0 17920 0 1 12544
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1491_
timestamp 1698431365
transform -1 0 18704 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1492_
timestamp 1698431365
transform 1 0 18592 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1493_
timestamp 1698431365
transform 1 0 18256 0 -1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1494_
timestamp 1698431365
transform 1 0 17248 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1495_
timestamp 1698431365
transform 1 0 15008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1496_
timestamp 1698431365
transform 1 0 17248 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1497_
timestamp 1698431365
transform -1 0 17136 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1498_
timestamp 1698431365
transform -1 0 19376 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1499_
timestamp 1698431365
transform 1 0 15680 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1500_
timestamp 1698431365
transform -1 0 11984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1501_
timestamp 1698431365
transform -1 0 15792 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1502_
timestamp 1698431365
transform 1 0 14336 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1503_
timestamp 1698431365
transform 1 0 12656 0 -1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1504_
timestamp 1698431365
transform 1 0 9744 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1505_
timestamp 1698431365
transform -1 0 5600 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1506_
timestamp 1698431365
transform -1 0 5264 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1507_
timestamp 1698431365
transform 1 0 9632 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1508_
timestamp 1698431365
transform -1 0 11088 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _1509_
timestamp 1698431365
transform 1 0 5936 0 -1 20384
box -86 -86 1766 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1510_
timestamp 1698431365
transform -1 0 7056 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1511_
timestamp 1698431365
transform -1 0 6384 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1512_
timestamp 1698431365
transform -1 0 3024 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1513_
timestamp 1698431365
transform 1 0 4592 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1514_
timestamp 1698431365
transform -1 0 6048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1515_
timestamp 1698431365
transform -1 0 6496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1516_
timestamp 1698431365
transform -1 0 8064 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1517_
timestamp 1698431365
transform -1 0 6608 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1518_
timestamp 1698431365
transform 1 0 4368 0 -1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1519_
timestamp 1698431365
transform 1 0 5488 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1520_
timestamp 1698431365
transform -1 0 15904 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1521_
timestamp 1698431365
transform 1 0 7616 0 1 23520
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1522_
timestamp 1698431365
transform 1 0 8288 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1523_
timestamp 1698431365
transform -1 0 9520 0 1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1524_
timestamp 1698431365
transform 1 0 7168 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1525_
timestamp 1698431365
transform 1 0 8288 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1526_
timestamp 1698431365
transform 1 0 9856 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _1527_
timestamp 1698431365
transform -1 0 9632 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1528_
timestamp 1698431365
transform -1 0 8288 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1529_
timestamp 1698431365
transform 1 0 9408 0 -1 23520
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1530_
timestamp 1698431365
transform 1 0 9856 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1531_
timestamp 1698431365
transform 1 0 7056 0 -1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1532_
timestamp 1698431365
transform -1 0 7616 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1533_
timestamp 1698431365
transform -1 0 6496 0 -1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1534_
timestamp 1698431365
transform 1 0 7840 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1535_
timestamp 1698431365
transform 1 0 6160 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1536_
timestamp 1698431365
transform -1 0 5936 0 -1 28224
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1537_
timestamp 1698431365
transform -1 0 7280 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or3_1  _1538_
timestamp 1698431365
transform -1 0 6608 0 1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1539_
timestamp 1698431365
transform 1 0 5152 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1540_
timestamp 1698431365
transform 1 0 4480 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1541_
timestamp 1698431365
transform -1 0 6384 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1542_
timestamp 1698431365
transform 1 0 4816 0 -1 29792
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1543_
timestamp 1698431365
transform -1 0 3024 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1544_
timestamp 1698431365
transform -1 0 7280 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1545_
timestamp 1698431365
transform -1 0 6608 0 1 31360
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1546_
timestamp 1698431365
transform 1 0 7728 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1547_
timestamp 1698431365
transform 1 0 5712 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1548_
timestamp 1698431365
transform 1 0 6160 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1549_
timestamp 1698431365
transform 1 0 5488 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1550_
timestamp 1698431365
transform -1 0 6832 0 -1 32928
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1551_
timestamp 1698431365
transform 1 0 5152 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1552_
timestamp 1698431365
transform -1 0 5824 0 -1 36064
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1553_
timestamp 1698431365
transform -1 0 5264 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1554_
timestamp 1698431365
transform -1 0 5600 0 -1 34496
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1555_
timestamp 1698431365
transform -1 0 8064 0 -1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1556_
timestamp 1698431365
transform 1 0 5488 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1557_
timestamp 1698431365
transform 1 0 6720 0 -1 29792
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _1558_
timestamp 1698431365
transform 1 0 7504 0 -1 29792
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _1559_
timestamp 1698431365
transform 1 0 6832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1560_
timestamp 1698431365
transform -1 0 7728 0 -1 39200
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1561_
timestamp 1698431365
transform 1 0 5600 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1562_
timestamp 1698431365
transform -1 0 6272 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1563_
timestamp 1698431365
transform 1 0 5712 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1564_
timestamp 1698431365
transform -1 0 5264 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1565_
timestamp 1698431365
transform 1 0 4816 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1566_
timestamp 1698431365
transform -1 0 8512 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1567_
timestamp 1698431365
transform 1 0 6272 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1568_
timestamp 1698431365
transform 1 0 4816 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1569_
timestamp 1698431365
transform -1 0 6272 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1570_
timestamp 1698431365
transform -1 0 6160 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1571_
timestamp 1698431365
transform 1 0 7728 0 -1 39200
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1572_
timestamp 1698431365
transform -1 0 9184 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1573_
timestamp 1698431365
transform 1 0 9632 0 -1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1574_
timestamp 1698431365
transform -1 0 8960 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1575_
timestamp 1698431365
transform -1 0 8736 0 1 39200
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1576_
timestamp 1698431365
transform -1 0 9744 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1577_
timestamp 1698431365
transform 1 0 8960 0 1 36064
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1578_
timestamp 1698431365
transform 1 0 9408 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1579_
timestamp 1698431365
transform 1 0 9408 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _1580_
timestamp 1698431365
transform -1 0 40768 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1581_
timestamp 1698431365
transform 1 0 9968 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1582_
timestamp 1698431365
transform -1 0 14000 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1583_
timestamp 1698431365
transform 1 0 9408 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _1584_
timestamp 1698431365
transform 1 0 8064 0 -1 36064
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _1585_
timestamp 1698431365
transform -1 0 9968 0 1 34496
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1586_
timestamp 1698431365
transform -1 0 10192 0 1 31360
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1587_
timestamp 1698431365
transform -1 0 9520 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _1588_
timestamp 1698431365
transform 1 0 9184 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1589_
timestamp 1698431365
transform -1 0 10752 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1590_
timestamp 1698431365
transform 1 0 10976 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1591_
timestamp 1698431365
transform 1 0 9968 0 1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1592_
timestamp 1698431365
transform 1 0 9072 0 1 32928
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1593_
timestamp 1698431365
transform 1 0 9408 0 -1 32928
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1594_
timestamp 1698431365
transform 1 0 10528 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1595_
timestamp 1698431365
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1596_
timestamp 1698431365
transform -1 0 10864 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _1597_
timestamp 1698431365
transform 1 0 9408 0 -1 28224
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1598_
timestamp 1698431365
transform -1 0 10416 0 1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1599_
timestamp 1698431365
transform 1 0 10416 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _1600_
timestamp 1698431365
transform 1 0 10640 0 -1 28224
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1601_
timestamp 1698431365
transform 1 0 10304 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _1602_
timestamp 1698431365
transform -1 0 10416 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1603_
timestamp 1698431365
transform -1 0 11648 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1604_
timestamp 1698431365
transform 1 0 38192 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1605_
timestamp 1698431365
transform -1 0 39088 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1606_
timestamp 1698431365
transform 1 0 38416 0 -1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1607_
timestamp 1698431365
transform 1 0 38752 0 1 31360
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1608_
timestamp 1698431365
transform 1 0 39200 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _1609_
timestamp 1698431365
transform 1 0 3472 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1610_
timestamp 1698431365
transform 1 0 30464 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1611_
timestamp 1698431365
transform -1 0 29792 0 1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _1612_
timestamp 1698431365
transform -1 0 30240 0 1 4704
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1613_
timestamp 1698431365
transform -1 0 25760 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1614_
timestamp 1698431365
transform 1 0 27776 0 1 4704
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1615_
timestamp 1698431365
transform -1 0 26320 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1616_
timestamp 1698431365
transform -1 0 22512 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1617_
timestamp 1698431365
transform -1 0 23072 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1618_
timestamp 1698431365
transform -1 0 22960 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1619_
timestamp 1698431365
transform 1 0 21056 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1620_
timestamp 1698431365
transform -1 0 19376 0 1 4704
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1621_
timestamp 1698431365
transform -1 0 29568 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1622_
timestamp 1698431365
transform 1 0 19376 0 -1 6272
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1623_
timestamp 1698431365
transform -1 0 19376 0 -1 6272
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1624_
timestamp 1698431365
transform 1 0 19488 0 -1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1625_
timestamp 1698431365
transform 1 0 20496 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1626_
timestamp 1698431365
transform 1 0 19936 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1627_
timestamp 1698431365
transform -1 0 19936 0 1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _1628_
timestamp 1698431365
transform -1 0 22848 0 1 7840
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _1629_
timestamp 1698431365
transform 1 0 23184 0 -1 7840
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1630_
timestamp 1698431365
transform -1 0 9184 0 1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _1631_
timestamp 1698431365
transform 1 0 7728 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1632_
timestamp 1698431365
transform 1 0 8064 0 -1 7840
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1633_
timestamp 1698431365
transform 1 0 38640 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1634_
timestamp 1698431365
transform -1 0 39088 0 1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1635_
timestamp 1698431365
transform 1 0 38640 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1636_
timestamp 1698431365
transform 1 0 36848 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1637_
timestamp 1698431365
transform -1 0 37408 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1638_
timestamp 1698431365
transform -1 0 41440 0 1 37632
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1639_
timestamp 1698431365
transform 1 0 36848 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1640_
timestamp 1698431365
transform -1 0 37968 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1641_
timestamp 1698431365
transform 1 0 36064 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1642_
timestamp 1698431365
transform 1 0 36848 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _1643_
timestamp 1698431365
transform 1 0 43344 0 1 42336
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1644_
timestamp 1698431365
transform 1 0 45248 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _1645_
timestamp 1698431365
transform 1 0 41888 0 -1 40768
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1646_
timestamp 1698431365
transform 1 0 43792 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1647_
timestamp 1698431365
transform -1 0 46032 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1648_
timestamp 1698431365
transform 1 0 44688 0 1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1649_
timestamp 1698431365
transform 1 0 43904 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1650_
timestamp 1698431365
transform 1 0 44688 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1651_
timestamp 1698431365
transform 1 0 45808 0 -1 43904
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1652_
timestamp 1698431365
transform 1 0 45920 0 1 39200
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1653_
timestamp 1698431365
transform 1 0 46592 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1654_
timestamp 1698431365
transform -1 0 43568 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1655_
timestamp 1698431365
transform -1 0 44352 0 -1 37632
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1656_
timestamp 1698431365
transform -1 0 43792 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1657_
timestamp 1698431365
transform 1 0 39760 0 -1 42336
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _1658_
timestamp 1698431365
transform 1 0 39872 0 -1 40768
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _1659_
timestamp 1698431365
transform 1 0 40768 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1660_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 44912 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1661_
timestamp 1698431365
transform 1 0 47824 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1662_
timestamp 1698431365
transform 1 0 50176 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1663_
timestamp 1698431365
transform 1 0 50176 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1664_
timestamp 1698431365
transform 1 0 50176 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1665_
timestamp 1698431365
transform 1 0 50176 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1666_
timestamp 1698431365
transform 1 0 50176 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1667_
timestamp 1698431365
transform -1 0 49952 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1668_
timestamp 1698431365
transform 1 0 50176 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1669_
timestamp 1698431365
transform 1 0 50176 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1670_
timestamp 1698431365
transform 1 0 50176 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1671_
timestamp 1698431365
transform 1 0 44016 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1672_
timestamp 1698431365
transform 1 0 40768 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1673_ $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 32928 0 -1 4704
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1674_
timestamp 1698431365
transform 1 0 41440 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1675_
timestamp 1698431365
transform -1 0 47936 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1676_
timestamp 1698431365
transform 1 0 42000 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1677_
timestamp 1698431365
transform 1 0 36960 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1678_
timestamp 1698431365
transform -1 0 36176 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1679_
timestamp 1698431365
transform 1 0 26992 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1680_
timestamp 1698431365
transform 1 0 29008 0 -1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1681_
timestamp 1698431365
transform 1 0 31472 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1682_
timestamp 1698431365
transform -1 0 40544 0 -1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1683_
timestamp 1698431365
transform 1 0 32704 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1684_
timestamp 1698431365
transform 1 0 26768 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1685_
timestamp 1698431365
transform 1 0 25536 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1686_
timestamp 1698431365
transform 1 0 21280 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1687_
timestamp 1698431365
transform 1 0 21280 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1688_
timestamp 1698431365
transform 1 0 19712 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1689_
timestamp 1698431365
transform 1 0 22512 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1690_
timestamp 1698431365
transform 1 0 23072 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1691_
timestamp 1698431365
transform 1 0 36736 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1692_
timestamp 1698431365
transform 1 0 35056 0 -1 32928
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1693_
timestamp 1698431365
transform 1 0 32928 0 -1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1694_
timestamp 1698431365
transform 1 0 29008 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1695_
timestamp 1698431365
transform 1 0 30016 0 1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1696_
timestamp 1698431365
transform 1 0 29232 0 -1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1697_
timestamp 1698431365
transform -1 0 29344 0 -1 29792
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1698_
timestamp 1698431365
transform -1 0 29008 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1699_
timestamp 1698431365
transform 1 0 30912 0 1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1700_
timestamp 1698431365
transform -1 0 51856 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1701_
timestamp 1698431365
transform 1 0 50176 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1702_
timestamp 1698431365
transform 1 0 45136 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1703_
timestamp 1698431365
transform 1 0 45920 0 1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1704_
timestamp 1698431365
transform 1 0 50176 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1705_
timestamp 1698431365
transform 1 0 50176 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1706_
timestamp 1698431365
transform 1 0 50176 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1707_
timestamp 1698431365
transform 1 0 50176 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1708_
timestamp 1698431365
transform 1 0 50176 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1709_
timestamp 1698431365
transform 1 0 45248 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1710_
timestamp 1698431365
transform 1 0 50176 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1711_
timestamp 1698431365
transform 1 0 50176 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1712_
timestamp 1698431365
transform 1 0 50176 0 -1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1713_
timestamp 1698431365
transform 1 0 44016 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1714_
timestamp 1698431365
transform 1 0 25312 0 1 31360
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1715_
timestamp 1698431365
transform 1 0 25200 0 1 34496
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1716_
timestamp 1698431365
transform 1 0 21504 0 1 36064
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1717_
timestamp 1698431365
transform 1 0 20272 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1718_
timestamp 1698431365
transform 1 0 19488 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1719_
timestamp 1698431365
transform 1 0 18816 0 -1 26656
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1720_
timestamp 1698431365
transform -1 0 20944 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1721_
timestamp 1698431365
transform 1 0 21504 0 1 23520
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1722_
timestamp 1698431365
transform 1 0 35056 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1723_
timestamp 1698431365
transform 1 0 33600 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1724_
timestamp 1698431365
transform 1 0 35168 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1725_
timestamp 1698431365
transform 1 0 29792 0 1 17248
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1726_
timestamp 1698431365
transform 1 0 26656 0 -1 15680
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1727_
timestamp 1698431365
transform 1 0 26320 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1728_
timestamp 1698431365
transform 1 0 30800 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1729_
timestamp 1698431365
transform 1 0 26096 0 -1 18816
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1730_
timestamp 1698431365
transform 1 0 28896 0 -1 42336
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1731_
timestamp 1698431365
transform 1 0 18816 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1732_
timestamp 1698431365
transform 1 0 25648 0 -1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1733_
timestamp 1698431365
transform 1 0 21392 0 -1 39200
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1734_
timestamp 1698431365
transform 1 0 19824 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1735_
timestamp 1698431365
transform -1 0 34160 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1736_
timestamp 1698431365
transform 1 0 29008 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1737_
timestamp 1698431365
transform 1 0 27664 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1738_
timestamp 1698431365
transform 1 0 32256 0 1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1739_
timestamp 1698431365
transform 1 0 15456 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1740_
timestamp 1698431365
transform 1 0 15680 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1741_
timestamp 1698431365
transform 1 0 16128 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1742_
timestamp 1698431365
transform 1 0 8512 0 1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1743_
timestamp 1698431365
transform 1 0 13328 0 1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1744_
timestamp 1698431365
transform 1 0 8736 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1745_
timestamp 1698431365
transform 1 0 13328 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1746_
timestamp 1698431365
transform 1 0 37296 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1747_
timestamp 1698431365
transform 1 0 33824 0 -1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1748_
timestamp 1698431365
transform -1 0 44352 0 1 50176
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1749_
timestamp 1698431365
transform 1 0 42672 0 -1 48608
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1750_
timestamp 1698431365
transform -1 0 47488 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1751_
timestamp 1698431365
transform 1 0 43568 0 -1 45472
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1752_
timestamp 1698431365
transform 1 0 40096 0 1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1753_
timestamp 1698431365
transform 1 0 35280 0 -1 47040
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1754_
timestamp 1698431365
transform 1 0 29008 0 1 43904
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1755_
timestamp 1698431365
transform 1 0 1568 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1756_
timestamp 1698431365
transform 1 0 1568 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1757_
timestamp 1698431365
transform 1 0 1568 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1758_
timestamp 1698431365
transform 1 0 1568 0 -1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1759_
timestamp 1698431365
transform 1 0 3808 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1760_
timestamp 1698431365
transform 1 0 6832 0 1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1761_
timestamp 1698431365
transform 1 0 9744 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1762_
timestamp 1698431365
transform 1 0 11200 0 -1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1763_
timestamp 1698431365
transform 1 0 13440 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1764_
timestamp 1698431365
transform 1 0 16800 0 1 10976
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1765_
timestamp 1698431365
transform 1 0 18368 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1766_
timestamp 1698431365
transform 1 0 15568 0 1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1767_
timestamp 1698431365
transform 1 0 11648 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1768_
timestamp 1698431365
transform 1 0 9408 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1769_
timestamp 1698431365
transform 1 0 1568 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1770_
timestamp 1698431365
transform 1 0 1568 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1771_
timestamp 1698431365
transform 1 0 12544 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1772_
timestamp 1698431365
transform 1 0 10304 0 -1 21952
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1773_
timestamp 1698431365
transform 1 0 1568 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1774_
timestamp 1698431365
transform 1 0 1568 0 -1 29792
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1775_
timestamp 1698431365
transform 1 0 1568 0 -1 32928
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1776_
timestamp 1698431365
transform 1 0 1568 0 1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1777_
timestamp 1698431365
transform 1 0 1568 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1778_
timestamp 1698431365
transform 1 0 4816 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1779_
timestamp 1698431365
transform 1 0 9744 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1780_
timestamp 1698431365
transform 1 0 10864 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1781_
timestamp 1698431365
transform 1 0 11088 0 -1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1782_
timestamp 1698431365
transform 1 0 10304 0 -1 34496
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1783_
timestamp 1698431365
transform 1 0 11760 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1784_
timestamp 1698431365
transform 1 0 10976 0 -1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1785_
timestamp 1698431365
transform 1 0 44688 0 1 31360
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1786_
timestamp 1698431365
transform 1 0 15456 0 1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1787_
timestamp 1698431365
transform 1 0 29120 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1788_
timestamp 1698431365
transform 1 0 25088 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1789_
timestamp 1698431365
transform 1 0 21392 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1790_
timestamp 1698431365
transform 1 0 17248 0 -1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1791_
timestamp 1698431365
transform 1 0 14336 0 1 4704
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1792_
timestamp 1698431365
transform 1 0 15232 0 1 6272
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1793_
timestamp 1698431365
transform 1 0 17248 0 -1 9408
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1794_
timestamp 1698431365
transform 1 0 22848 0 1 7840
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _1795_
timestamp 1698431365
transform 1 0 7616 0 1 6272
box -86 -86 3558 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1796_
timestamp 1698431365
transform 1 0 37296 0 -1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1797_
timestamp 1698431365
transform 1 0 33376 0 1 40768
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1798_
timestamp 1698431365
transform 1 0 33376 0 1 37632
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1799_
timestamp 1698431365
transform -1 0 48384 0 -1 42336
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1800_
timestamp 1698431365
transform -1 0 45920 0 -1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1801_
timestamp 1698431365
transform -1 0 49840 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1802_
timestamp 1698431365
transform -1 0 45472 0 -1 36064
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _1803_
timestamp 1698431365
transform -1 0 41552 0 1 39200
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0830__I $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 40992 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0831__I
timestamp 1698431365
transform 1 0 40208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0836__I
timestamp 1698431365
transform 1 0 33152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__A1
timestamp 1698431365
transform 1 0 33936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0838__B2
timestamp 1698431365
transform -1 0 34832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0842__A1
timestamp 1698431365
transform 1 0 37072 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0844__B2
timestamp 1698431365
transform 1 0 34832 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0848__A1
timestamp 1698431365
transform -1 0 39088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0856__I
timestamp 1698431365
transform 1 0 46928 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0857__I
timestamp 1698431365
transform 1 0 44016 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0859__A2
timestamp 1698431365
transform 1 0 43904 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A1
timestamp 1698431365
transform 1 0 44912 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0860__A2
timestamp 1698431365
transform 1 0 45360 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0861__A2
timestamp 1698431365
transform 1 0 42112 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0862__I
timestamp 1698431365
transform 1 0 45360 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0864__A1
timestamp 1698431365
transform -1 0 45472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0866__A1
timestamp 1698431365
transform -1 0 45584 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0867__I
timestamp 1698431365
transform -1 0 39760 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0868__I
timestamp 1698431365
transform -1 0 40768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0871__A2
timestamp 1698431365
transform 1 0 42112 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0873__A2
timestamp 1698431365
transform 1 0 49056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0874__I
timestamp 1698431365
transform 1 0 47376 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0875__A1
timestamp 1698431365
transform 1 0 49952 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0879__A1
timestamp 1698431365
transform -1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0880__I
timestamp 1698431365
transform 1 0 41664 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0881__I
timestamp 1698431365
transform 1 0 41664 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0882__I
timestamp 1698431365
transform 1 0 45920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0883__A2
timestamp 1698431365
transform 1 0 50624 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0888__A2
timestamp 1698431365
transform 1 0 50400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0902__I
timestamp 1698431365
transform 1 0 46368 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0907__I
timestamp 1698431365
transform 1 0 45584 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0914__A1
timestamp 1698431365
transform 1 0 48832 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0921__A3
timestamp 1698431365
transform 1 0 44240 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0923__I
timestamp 1698431365
transform -1 0 37744 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0924__C
timestamp 1698431365
transform -1 0 49056 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0930__C
timestamp 1698431365
transform 1 0 47712 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0936__C
timestamp 1698431365
transform -1 0 49280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0940__C
timestamp 1698431365
transform 1 0 44016 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0942__I
timestamp 1698431365
transform 1 0 40544 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0947__A2
timestamp 1698431365
transform 1 0 42448 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0951__A1
timestamp 1698431365
transform -1 0 43456 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0952__I
timestamp 1698431365
transform 1 0 23968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0954__I
timestamp 1698431365
transform 1 0 26432 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__A1
timestamp 1698431365
transform 1 0 37184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0956__A2
timestamp 1698431365
transform -1 0 36960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0959__A2
timestamp 1698431365
transform 1 0 43232 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0964__C
timestamp 1698431365
transform 1 0 40768 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0966__A2
timestamp 1698431365
transform 1 0 46816 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0971__B
timestamp 1698431365
transform -1 0 43344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0975__C
timestamp 1698431365
transform 1 0 41216 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__0988__B
timestamp 1698431365
transform -1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__A1
timestamp 1698431365
transform 1 0 38752 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1002__B
timestamp 1698431365
transform 1 0 39200 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1003__A3
timestamp 1698431365
transform 1 0 46592 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1006__A1
timestamp 1698431365
transform -1 0 35952 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1007__C
timestamp 1698431365
transform 1 0 33152 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1009__I
timestamp 1698431365
transform 1 0 26544 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1011__A1
timestamp 1698431365
transform 1 0 27888 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1016__I
timestamp 1698431365
transform 1 0 25984 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1018__A1
timestamp 1698431365
transform 1 0 24752 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1019__I
timestamp 1698431365
transform 1 0 22288 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1023__A1
timestamp 1698431365
transform 1 0 24640 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1034__B
timestamp 1698431365
transform -1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__A1
timestamp 1698431365
transform 1 0 39872 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1035__B
timestamp 1698431365
transform 1 0 39424 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1036__I0
timestamp 1698431365
transform -1 0 39872 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1038__I
timestamp 1698431365
transform 1 0 26880 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A1
timestamp 1698431365
transform 1 0 44912 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1039__A2
timestamp 1698431365
transform -1 0 45584 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1040__I
timestamp 1698431365
transform 1 0 44464 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1042__A1
timestamp 1698431365
transform -1 0 36512 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1044__A1
timestamp 1698431365
transform 1 0 35168 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1046__A1
timestamp 1698431365
transform 1 0 33712 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1048__I
timestamp 1698431365
transform -1 0 26768 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1051__A1
timestamp 1698431365
transform 1 0 31920 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1052__A1
timestamp 1698431365
transform 1 0 34272 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1055__A1
timestamp 1698431365
transform 1 0 31472 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1056__A1
timestamp 1698431365
transform 1 0 29904 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1059__A1
timestamp 1698431365
transform 1 0 31920 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1060__A1
timestamp 1698431365
transform 1 0 30912 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1063__A1
timestamp 1698431365
transform -1 0 31920 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1065__A1
timestamp 1698431365
transform 1 0 29344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1069__A1
timestamp 1698431365
transform 1 0 30240 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1070__A1
timestamp 1698431365
transform 1 0 30912 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1073__A1
timestamp 1698431365
transform -1 0 30464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1074__A1
timestamp 1698431365
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1076__I
timestamp 1698431365
transform 1 0 47152 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1077__A1
timestamp 1698431365
transform -1 0 31808 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1078__A1
timestamp 1698431365
transform -1 0 31584 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1080__A2
timestamp 1698431365
transform 1 0 46480 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1081__I
timestamp 1698431365
transform -1 0 47712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1082__I
timestamp 1698431365
transform -1 0 41664 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1083__I
timestamp 1698431365
transform 1 0 49056 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1084__I
timestamp 1698431365
transform 1 0 44464 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1087__I
timestamp 1698431365
transform 1 0 42224 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1090__A1
timestamp 1698431365
transform 1 0 38080 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1091__A2
timestamp 1698431365
transform -1 0 43456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1093__I
timestamp 1698431365
transform -1 0 26320 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__B1
timestamp 1698431365
transform 1 0 37520 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1094__B2
timestamp 1698431365
transform 1 0 37072 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1097__I
timestamp 1698431365
transform 1 0 41664 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1099__I
timestamp 1698431365
transform 1 0 26768 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1100__A1
timestamp 1698431365
transform 1 0 44240 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1102__A2
timestamp 1698431365
transform 1 0 44016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__A1
timestamp 1698431365
transform 1 0 36624 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1104__B2
timestamp 1698431365
transform -1 0 37296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__A1
timestamp 1698431365
transform 1 0 35728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__B1
timestamp 1698431365
transform 1 0 36624 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1109__B2
timestamp 1698431365
transform 1 0 36176 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1112__A1
timestamp 1698431365
transform -1 0 37520 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1114__B2
timestamp 1698431365
transform 1 0 37744 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1115__B
timestamp 1698431365
transform 1 0 48384 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__A1
timestamp 1698431365
transform 1 0 35728 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__B1
timestamp 1698431365
transform -1 0 37296 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1117__B2
timestamp 1698431365
transform 1 0 36176 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1122__B
timestamp 1698431365
transform 1 0 48160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1126__I
timestamp 1698431365
transform -1 0 23968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__A1
timestamp 1698431365
transform 1 0 25088 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1127__B1
timestamp 1698431365
transform 1 0 24640 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__A1
timestamp 1698431365
transform -1 0 35840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1128__B2
timestamp 1698431365
transform 1 0 35168 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1129__A3
timestamp 1698431365
transform -1 0 42896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1133__I
timestamp 1698431365
transform 1 0 25312 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1134__A1
timestamp 1698431365
transform -1 0 24640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__A1
timestamp 1698431365
transform 1 0 37184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1136__B2
timestamp 1698431365
transform 1 0 37632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1137__A3
timestamp 1698431365
transform 1 0 42560 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1141__B2
timestamp 1698431365
transform 1 0 21840 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1142__A1
timestamp 1698431365
transform -1 0 34160 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1143__A3
timestamp 1698431365
transform -1 0 42448 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1146__I
timestamp 1698431365
transform 1 0 48160 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1148__B2
timestamp 1698431365
transform 1 0 22960 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1149__A1
timestamp 1698431365
transform -1 0 34496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1150__A3
timestamp 1698431365
transform 1 0 41328 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1151__B
timestamp 1698431365
transform -1 0 48496 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1152__A1
timestamp 1698431365
transform 1 0 49280 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1154__B2
timestamp 1698431365
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__A1
timestamp 1698431365
transform -1 0 35392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1155__B2
timestamp 1698431365
transform 1 0 35392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1157__B
timestamp 1698431365
transform -1 0 50288 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1158__A1
timestamp 1698431365
transform 1 0 52080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1160__A2
timestamp 1698431365
transform -1 0 16576 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1161__A2
timestamp 1698431365
transform 1 0 20160 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1163__A2
timestamp 1698431365
transform -1 0 20160 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1165__A2
timestamp 1698431365
transform 1 0 17920 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1166__A2
timestamp 1698431365
transform 1 0 21392 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1168__A2
timestamp 1698431365
transform -1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1171__A2
timestamp 1698431365
transform -1 0 33376 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1172__A2
timestamp 1698431365
transform 1 0 32928 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1173__A2
timestamp 1698431365
transform -1 0 29344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1174__A2
timestamp 1698431365
transform 1 0 30016 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1176__A2
timestamp 1698431365
transform 1 0 29232 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1177__A2
timestamp 1698431365
transform -1 0 26880 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1178__A2
timestamp 1698431365
transform 1 0 29232 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1179__A2
timestamp 1698431365
transform 1 0 26880 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1182__A2
timestamp 1698431365
transform 1 0 32256 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1183__A2
timestamp 1698431365
transform 1 0 48160 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1185__I
timestamp 1698431365
transform -1 0 37184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1187__A2
timestamp 1698431365
transform 1 0 46368 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1188__B
timestamp 1698431365
transform 1 0 46144 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1191__A1
timestamp 1698431365
transform -1 0 51744 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1193__A3
timestamp 1698431365
transform -1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1194__B
timestamp 1698431365
transform 1 0 49728 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1199__A1
timestamp 1698431365
transform 1 0 47488 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1201__A1
timestamp 1698431365
transform -1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1203__I
timestamp 1698431365
transform 1 0 26880 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__A1
timestamp 1698431365
transform 1 0 37856 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1206__C
timestamp 1698431365
transform 1 0 39200 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A1
timestamp 1698431365
transform 1 0 27328 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1207__A2
timestamp 1698431365
transform 1 0 26208 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1209__A1
timestamp 1698431365
transform 1 0 26208 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1210__I
timestamp 1698431365
transform 1 0 20384 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__A1
timestamp 1698431365
transform 1 0 26432 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1212__C
timestamp 1698431365
transform 1 0 24640 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1213__A1
timestamp 1698431365
transform -1 0 26432 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1214__A2
timestamp 1698431365
transform 1 0 25760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1216__A1
timestamp 1698431365
transform 1 0 24192 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1217__B
timestamp 1698431365
transform 1 0 24640 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1218__A1
timestamp 1698431365
transform -1 0 24192 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1219__A1
timestamp 1698431365
transform 1 0 21840 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1220__B
timestamp 1698431365
transform 1 0 23744 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1221__A1
timestamp 1698431365
transform 1 0 23520 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1226__A1
timestamp 1698431365
transform 1 0 21392 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1229__A1
timestamp 1698431365
transform -1 0 19040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1230__A1
timestamp 1698431365
transform 1 0 19152 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1232__A1
timestamp 1698431365
transform 1 0 21056 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1233__A1
timestamp 1698431365
transform 1 0 20272 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1235__A1
timestamp 1698431365
transform 1 0 23408 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1236__A1
timestamp 1698431365
transform 1 0 21840 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1243__A1
timestamp 1698431365
transform -1 0 34944 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1246__A1
timestamp 1698431365
transform -1 0 33040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1249__A1
timestamp 1698431365
transform 1 0 33936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1252__A1
timestamp 1698431365
transform 1 0 32144 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1254__A1
timestamp 1698431365
transform 1 0 27664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1255__A1
timestamp 1698431365
transform 1 0 30016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1257__A1
timestamp 1698431365
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__A1
timestamp 1698431365
transform 1 0 34720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1260__B
timestamp 1698431365
transform 1 0 35168 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1262__A1
timestamp 1698431365
transform 1 0 29232 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1263__A1
timestamp 1698431365
transform 1 0 29792 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1267__I
timestamp 1698431365
transform 1 0 27888 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1268__I
timestamp 1698431365
transform 1 0 34832 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1271__I
timestamp 1698431365
transform 1 0 24528 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1274__A1
timestamp 1698431365
transform 1 0 30464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1282__I
timestamp 1698431365
transform 1 0 21616 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1283__I
timestamp 1698431365
transform 1 0 20720 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1286__I
timestamp 1698431365
transform 1 0 16800 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1289__A2
timestamp 1698431365
transform 1 0 22960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1291__A1
timestamp 1698431365
transform 1 0 27328 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1293__A2
timestamp 1698431365
transform -1 0 24080 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1299__C
timestamp 1698431365
transform 1 0 22624 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1302__A2
timestamp 1698431365
transform 1 0 38640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1303__B
timestamp 1698431365
transform 1 0 26208 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1305__I
timestamp 1698431365
transform 1 0 25424 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1308__I
timestamp 1698431365
transform 1 0 40992 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1314__B
timestamp 1698431365
transform 1 0 27552 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1328__B
timestamp 1698431365
transform 1 0 23072 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1335__I
timestamp 1698431365
transform -1 0 11648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1340__B
timestamp 1698431365
transform -1 0 19824 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1341__A1
timestamp 1698431365
transform 1 0 18032 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1344__A1
timestamp 1698431365
transform -1 0 19936 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1349__B
timestamp 1698431365
transform 1 0 15344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1351__A1
timestamp 1698431365
transform 1 0 13552 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1353__A1
timestamp 1698431365
transform 1 0 12768 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1366__B
timestamp 1698431365
transform -1 0 16128 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1367__C
timestamp 1698431365
transform 1 0 15568 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1370__A1
timestamp 1698431365
transform 1 0 38528 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1378__I
timestamp 1698431365
transform 1 0 41776 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1390__A1
timestamp 1698431365
transform 1 0 40544 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1391__B
timestamp 1698431365
transform 1 0 39648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1393__A2
timestamp 1698431365
transform 1 0 32704 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1396__A1
timestamp 1698431365
transform 1 0 28560 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1398__A2
timestamp 1698431365
transform 1 0 17472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1399__A2
timestamp 1698431365
transform -1 0 19376 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1401__A2
timestamp 1698431365
transform 1 0 16688 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1403__A2
timestamp 1698431365
transform 1 0 18816 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1404__A2
timestamp 1698431365
transform -1 0 17248 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1405__A2
timestamp 1698431365
transform 1 0 17808 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1406__A2
timestamp 1698431365
transform 1 0 15904 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1410__A2
timestamp 1698431365
transform 1 0 19376 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__A1
timestamp 1698431365
transform -1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1411__A2
timestamp 1698431365
transform 1 0 19936 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A1
timestamp 1698431365
transform 1 0 16800 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1412__A2
timestamp 1698431365
transform 1 0 18704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1415__A2
timestamp 1698431365
transform 1 0 15456 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1416__A2
timestamp 1698431365
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1417__A2
timestamp 1698431365
transform 1 0 15456 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A1
timestamp 1698431365
transform 1 0 12992 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1418__A2
timestamp 1698431365
transform 1 0 14560 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1421__I
timestamp 1698431365
transform 1 0 8960 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1423__A1
timestamp 1698431365
transform 1 0 41664 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1425__A2
timestamp 1698431365
transform 1 0 9632 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1431__A1
timestamp 1698431365
transform 1 0 15008 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1433__A2
timestamp 1698431365
transform 1 0 8512 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1435__A2
timestamp 1698431365
transform 1 0 8512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1439__I
timestamp 1698431365
transform -1 0 15008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1445__I
timestamp 1698431365
transform 1 0 31136 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1446__C
timestamp 1698431365
transform 1 0 7280 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1449__I
timestamp 1698431365
transform 1 0 10304 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1451__B
timestamp 1698431365
transform -1 0 7728 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1454__A2
timestamp 1698431365
transform 1 0 11984 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1457__C
timestamp 1698431365
transform 1 0 6944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1462__I
timestamp 1698431365
transform 1 0 8736 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1463__B
timestamp 1698431365
transform 1 0 7840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A1
timestamp 1698431365
transform 1 0 11872 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1466__A2
timestamp 1698431365
transform -1 0 11648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1468__C
timestamp 1698431365
transform -1 0 12096 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1470__I
timestamp 1698431365
transform 1 0 16576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1472__A1
timestamp 1698431365
transform -1 0 13552 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1473__C
timestamp 1698431365
transform 1 0 13216 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1477__A1
timestamp 1698431365
transform 1 0 15120 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1483__A1
timestamp 1698431365
transform -1 0 17696 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1489__A1
timestamp 1698431365
transform -1 0 20384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1493__A1
timestamp 1698431365
transform -1 0 19824 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1497__A1
timestamp 1698431365
transform 1 0 18144 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1502__A1
timestamp 1698431365
transform 1 0 15680 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1505__I
timestamp 1698431365
transform 1 0 4704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1512__A1
timestamp 1698431365
transform 1 0 3248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1513__I
timestamp 1698431365
transform 1 0 5264 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1519__B
timestamp 1698431365
transform 1 0 6608 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1521__A3
timestamp 1698431365
transform 1 0 7392 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1525__A1
timestamp 1698431365
transform 1 0 9184 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1526__I
timestamp 1698431365
transform 1 0 9632 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A1
timestamp 1698431365
transform 1 0 9856 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A3
timestamp 1698431365
transform 1 0 7168 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1527__A4
timestamp 1698431365
transform 1 0 7616 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1529__A1
timestamp 1698431365
transform 1 0 11312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1534__A1
timestamp 1698431365
transform 1 0 8624 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1539__B
timestamp 1698431365
transform 1 0 6272 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1543__A1
timestamp 1698431365
transform 1 0 3248 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1551__B
timestamp 1698431365
transform 1 0 7056 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1555__I
timestamp 1698431365
transform 1 0 8064 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1581__B
timestamp 1698431365
transform 1 0 10864 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1590__A1
timestamp 1698431365
transform 1 0 11872 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1594__B
timestamp 1698431365
transform 1 0 11648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1600__C
timestamp 1698431365
transform 1 0 11760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1603__C
timestamp 1698431365
transform 1 0 11872 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1606__A1
timestamp 1698431365
transform 1 0 38192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1608__B
timestamp 1698431365
transform -1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1610__A1
timestamp 1698431365
transform -1 0 31584 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__A1
timestamp 1698431365
transform 1 0 28784 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1612__C
timestamp 1698431365
transform -1 0 30688 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1631__A1
timestamp 1698431365
transform -1 0 9632 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1632__A1
timestamp 1698431365
transform -1 0 9072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1635__B
timestamp 1698431365
transform 1 0 39760 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1653__B
timestamp 1698431365
transform 1 0 46368 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1656__B
timestamp 1698431365
transform 1 0 42672 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1659__B
timestamp 1698431365
transform -1 0 41888 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1664__CLK
timestamp 1698431365
transform 1 0 49952 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1665__CLK
timestamp 1698431365
transform 1 0 49392 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1666__CLK
timestamp 1698431365
transform 1 0 49952 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1667__CLK
timestamp 1698431365
transform 1 0 50176 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1668__CLK
timestamp 1698431365
transform 1 0 49952 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1669__CLK
timestamp 1698431365
transform 1 0 49952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1670__CLK
timestamp 1698431365
transform 1 0 49504 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1671__CLK
timestamp 1698431365
transform 1 0 47488 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1672__CLK
timestamp 1698431365
transform 1 0 40544 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1673__CLK
timestamp 1698431365
transform 1 0 36400 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1674__CLK
timestamp 1698431365
transform 1 0 41216 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1675__CLK
timestamp 1698431365
transform 1 0 47936 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1676__CLK
timestamp 1698431365
transform 1 0 41776 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1677__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1678__CLK
timestamp 1698431365
transform 1 0 36176 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1679__CLK
timestamp 1698431365
transform 1 0 26768 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1680__CLK
timestamp 1698431365
transform 1 0 28784 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1681__CLK
timestamp 1698431365
transform 1 0 31248 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1682__CLK
timestamp 1698431365
transform 1 0 40992 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1683__CLK
timestamp 1698431365
transform 1 0 35952 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1684__CLK
timestamp 1698431365
transform 1 0 26544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1685__CLK
timestamp 1698431365
transform 1 0 25312 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1686__CLK
timestamp 1698431365
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1687__CLK
timestamp 1698431365
transform 1 0 24752 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1688__CLK
timestamp 1698431365
transform 1 0 23184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1689__CLK
timestamp 1698431365
transform 1 0 25984 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1690__CLK
timestamp 1698431365
transform 1 0 22288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1691__CLK
timestamp 1698431365
transform 1 0 40208 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1692__CLK
timestamp 1698431365
transform 1 0 38752 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1693__CLK
timestamp 1698431365
transform 1 0 36400 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1694__CLK
timestamp 1698431365
transform 1 0 32704 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1695__CLK
timestamp 1698431365
transform 1 0 33712 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1696__CLK
timestamp 1698431365
transform 1 0 33152 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1697__CLK
timestamp 1698431365
transform -1 0 29792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1698__CLK
timestamp 1698431365
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1699__CLK
timestamp 1698431365
transform 1 0 34720 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1700__CLK
timestamp 1698431365
transform 1 0 49056 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1707__CLK
timestamp 1698431365
transform 1 0 49952 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1709__CLK
timestamp 1698431365
transform 1 0 48720 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1710__CLK
timestamp 1698431365
transform 1 0 49952 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1711__CLK
timestamp 1698431365
transform 1 0 49952 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1712__CLK
timestamp 1698431365
transform 1 0 49952 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1714__CLK
timestamp 1698431365
transform 1 0 29232 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1715__CLK
timestamp 1698431365
transform 1 0 28672 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1720__CLK
timestamp 1698431365
transform 1 0 20944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1721__CLK
timestamp 1698431365
transform 1 0 25200 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1722__CLK
timestamp 1698431365
transform 1 0 38528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1723__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1724__CLK
timestamp 1698431365
transform 1 0 38864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1725__CLK
timestamp 1698431365
transform 1 0 29568 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1726__CLK
timestamp 1698431365
transform 1 0 26432 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1727__CLK
timestamp 1698431365
transform 1 0 26096 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1728__CLK
timestamp 1698431365
transform 1 0 30576 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1729__CLK
timestamp 1698431365
transform 1 0 25872 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1730__CLK
timestamp 1698431365
transform 1 0 32368 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1731__CLK
timestamp 1698431365
transform 1 0 18592 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1732__CLK
timestamp 1698431365
transform 1 0 29120 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1734__CLK
timestamp 1698431365
transform 1 0 19600 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1735__CLK
timestamp 1698431365
transform 1 0 34384 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1736__CLK
timestamp 1698431365
transform 1 0 32256 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1737__CLK
timestamp 1698431365
transform 1 0 30912 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1738__CLK
timestamp 1698431365
transform 1 0 35728 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1739__CLK
timestamp 1698431365
transform 1 0 18928 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1740__CLK
timestamp 1698431365
transform 1 0 19152 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1741__CLK
timestamp 1698431365
transform 1 0 19600 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1742__CLK
timestamp 1698431365
transform -1 0 11984 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1743__CLK
timestamp 1698431365
transform 1 0 16800 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1744__CLK
timestamp 1698431365
transform 1 0 12208 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1745__CLK
timestamp 1698431365
transform 1 0 16576 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1746__CLK
timestamp 1698431365
transform 1 0 37072 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1747__CLK
timestamp 1698431365
transform 1 0 37072 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1748__CLK
timestamp 1698431365
transform 1 0 44912 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1749__CLK
timestamp 1698431365
transform 1 0 46144 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1750__CLK
timestamp 1698431365
transform 1 0 47712 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1751__CLK
timestamp 1698431365
transform 1 0 47040 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1752__CLK
timestamp 1698431365
transform 1 0 44240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1753__CLK
timestamp 1698431365
transform 1 0 38528 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1754__CLK
timestamp 1698431365
transform 1 0 32480 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1755__CLK
timestamp 1698431365
transform 1 0 5040 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1756__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1757__CLK
timestamp 1698431365
transform 1 0 4816 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1758__CLK
timestamp 1698431365
transform 1 0 5040 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1759__CLK
timestamp 1698431365
transform 1 0 7728 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1760__CLK
timestamp 1698431365
transform 1 0 10304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1761__CLK
timestamp 1698431365
transform 1 0 13552 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1762__CLK
timestamp 1698431365
transform 1 0 14672 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1763__CLK
timestamp 1698431365
transform 1 0 16688 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1764__CLK
timestamp 1698431365
transform 1 0 16576 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1765__CLK
timestamp 1698431365
transform 1 0 21616 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1766__CLK
timestamp 1698431365
transform 1 0 15344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1767__CLK
timestamp 1698431365
transform 1 0 15120 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1768__CLK
timestamp 1698431365
transform 1 0 12656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1769__CLK
timestamp 1698431365
transform 1 0 5040 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1770__CLK
timestamp 1698431365
transform 1 0 5712 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1771__CLK
timestamp 1698431365
transform 1 0 12320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1772__CLK
timestamp 1698431365
transform 1 0 14000 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1773__CLK
timestamp 1698431365
transform 1 0 5040 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1774__CLK
timestamp 1698431365
transform -1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1775__CLK
timestamp 1698431365
transform 1 0 4816 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1776__CLK
timestamp 1698431365
transform 1 0 4816 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1777__CLK
timestamp 1698431365
transform 1 0 4816 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1778__CLK
timestamp 1698431365
transform 1 0 8288 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1779__CLK
timestamp 1698431365
transform 1 0 12992 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1780__CLK
timestamp 1698431365
transform 1 0 14336 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1781__CLK
timestamp 1698431365
transform 1 0 11088 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1782__CLK
timestamp 1698431365
transform 1 0 13776 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1783__CLK
timestamp 1698431365
transform 1 0 12208 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1784__CLK
timestamp 1698431365
transform 1 0 10080 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__CLK
timestamp 1698431365
transform -1 0 15680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1786__D
timestamp 1698431365
transform 1 0 15232 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1787__CLK
timestamp 1698431365
transform -1 0 29120 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1788__CLK
timestamp 1698431365
transform -1 0 25088 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1789__CLK
timestamp 1698431365
transform 1 0 24640 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1790__CLK
timestamp 1698431365
transform 1 0 16800 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1791__CLK
timestamp 1698431365
transform 1 0 17808 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1792__CLK
timestamp 1698431365
transform 1 0 15008 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1793__CLK
timestamp 1698431365
transform 1 0 17024 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1794__CLK
timestamp 1698431365
transform 1 0 26320 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1795__CLK
timestamp 1698431365
transform 1 0 11312 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1796__CLK
timestamp 1698431365
transform 1 0 37072 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1797__CLK
timestamp 1698431365
transform 1 0 36624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1798__CLK
timestamp 1698431365
transform 1 0 37968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1799__CLK
timestamp 1698431365
transform 1 0 48832 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__1803__CLK
timestamp 1698431365
transform 1 0 41776 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 26880 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_0_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_1_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 16464 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_2_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_3_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 25312 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_4_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 13440 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_5_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 12992 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_6_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 20272 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_7_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 19152 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_8_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 39200 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_9_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 37968 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_10_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 45360 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_11_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 45248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_12_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 34832 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_13_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 35392 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_14_0_wb_clk_i_I
timestamp 1698431365
transform -1 0 43792 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_4_15_0_wb_clk_i_I
timestamp 1698431365
transform 1 0 44240 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input1_I
timestamp 1698431365
transform -1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input2_I
timestamp 1698431365
transform -1 0 52528 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input3_I
timestamp 1698431365
transform -1 0 51408 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input4_I
timestamp 1698431365
transform -1 0 52752 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input5_I
timestamp 1698431365
transform -1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input6_I
timestamp 1698431365
transform -1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input7_I
timestamp 1698431365
transform -1 0 53424 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input8_I
timestamp 1698431365
transform -1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input9_I
timestamp 1698431365
transform -1 0 53424 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input10_I
timestamp 1698431365
transform -1 0 53424 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input11_I
timestamp 1698431365
transform -1 0 53424 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input12_I
timestamp 1698431365
transform 1 0 53200 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input13_I
timestamp 1698431365
transform -1 0 52752 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input14_I
timestamp 1698431365
transform -1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input15_I
timestamp 1698431365
transform -1 0 2800 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_input16_I
timestamp 1698431365
transform -1 0 41328 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output17_I
timestamp 1698431365
transform -1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output26_I
timestamp 1698431365
transform -1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output27_I
timestamp 1698431365
transform 1 0 14896 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 27104 0 -1 28224
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_0_0_wb_clk_i $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 16464 0 1 14112
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_1_0_wb_clk_i
timestamp 1698431365
transform 1 0 13328 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_2_0_wb_clk_i
timestamp 1698431365
transform -1 0 24864 0 -1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_3_0_wb_clk_i
timestamp 1698431365
transform -1 0 24864 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_4_0_wb_clk_i
timestamp 1698431365
transform -1 0 12544 0 -1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_5_0_wb_clk_i
timestamp 1698431365
transform -1 0 12992 0 1 29792
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_6_0_wb_clk_i
timestamp 1698431365
transform 1 0 17136 0 1 31360
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_7_0_wb_clk_i
timestamp 1698431365
transform -1 0 18368 0 1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_8_0_wb_clk_i
timestamp 1698431365
transform -1 0 42336 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_9_0_wb_clk_i
timestamp 1698431365
transform -1 0 41104 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_10_0_wb_clk_i
timestamp 1698431365
transform 1 0 45584 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_11_0_wb_clk_i
timestamp 1698431365
transform 1 0 45472 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_12_0_wb_clk_i
timestamp 1698431365
transform -1 0 37968 0 -1 39200
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_13_0_wb_clk_i
timestamp 1698431365
transform -1 0 38304 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_14_0_wb_clk_i
timestamp 1698431365
transform 1 0 44352 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_8  clkbuf_4_15_0_wb_clk_i
timestamp 1698431365
transform 1 0 44688 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_2 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1568 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_10 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 2464 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_19
timestamp 1698431365
transform 1 0 3472 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_27 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4368 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_31 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 4816 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_33
timestamp 1698431365
transform 1 0 5040 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_96
timestamp 1698431365
transform 1 0 12096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_100
timestamp 1698431365
transform 1 0 12544 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698431365
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_142 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 17248 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_158
timestamp 1698431365
transform 1 0 19040 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_166
timestamp 1698431365
transform 1 0 19936 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_172
timestamp 1698431365
transform 1 0 20608 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_177
timestamp 1698431365
transform 1 0 21168 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_193
timestamp 1698431365
transform 1 0 22960 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_201
timestamp 1698431365
transform 1 0 23856 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_203
timestamp 1698431365
transform 1 0 24080 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_206
timestamp 1698431365
transform 1 0 24416 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_212
timestamp 1698431365
transform 1 0 25088 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_217
timestamp 1698431365
transform 1 0 25648 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_233
timestamp 1698431365
transform 1 0 27440 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_237
timestamp 1698431365
transform 1 0 27888 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_240
timestamp 1698431365
transform 1 0 28224 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_244
timestamp 1698431365
transform 1 0 28672 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_248
timestamp 1698431365
transform 1 0 29120 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_252
timestamp 1698431365
transform 1 0 29568 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_257
timestamp 1698431365
transform 1 0 30128 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_265
timestamp 1698431365
transform 1 0 31024 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_269
timestamp 1698431365
transform 1 0 31472 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698431365
transform 1 0 31696 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_274
timestamp 1698431365
transform 1 0 32032 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_290
timestamp 1698431365
transform 1 0 33824 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_298
timestamp 1698431365
transform 1 0 34720 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_302
timestamp 1698431365
transform 1 0 35168 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_334
timestamp 1698431365
transform 1 0 38752 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_350
timestamp 1698431365
transform 1 0 40544 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_366
timestamp 1698431365
transform 1 0 42336 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_370
timestamp 1698431365
transform 1 0 42784 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_382
timestamp 1698431365
transform 1 0 44128 0 1 3136
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_398
timestamp 1698431365
transform 1 0 45920 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_444
timestamp 1698431365
transform 1 0 51072 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_452
timestamp 1698431365
transform 1 0 51968 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_454
timestamp 1698431365
transform 1 0 52192 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_2
timestamp 1698431365
transform 1 0 1568 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_18
timestamp 1698431365
transform 1 0 3360 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_23
timestamp 1698431365
transform 1 0 3920 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_55
timestamp 1698431365
transform 1 0 7504 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_63
timestamp 1698431365
transform 1 0 8400 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_67
timestamp 1698431365
transform 1 0 8848 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_69
timestamp 1698431365
transform 1 0 9072 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_72
timestamp 1698431365
transform 1 0 9408 0 -1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_88
timestamp 1698431365
transform 1 0 11200 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_92
timestamp 1698431365
transform 1 0 11648 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_119
timestamp 1698431365
transform 1 0 14672 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_123
timestamp 1698431365
transform 1 0 15120 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_131
timestamp 1698431365
transform 1 0 16016 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_135
timestamp 1698431365
transform 1 0 16464 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_137
timestamp 1698431365
transform 1 0 16688 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_171
timestamp 1698431365
transform 1 0 20496 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698431365
transform 1 0 24640 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_241
timestamp 1698431365
transform 1 0 28336 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_247
timestamp 1698431365
transform 1 0 29008 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_277
timestamp 1698431365
transform 1 0 32368 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_279
timestamp 1698431365
transform 1 0 32592 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_313
timestamp 1698431365
transform 1 0 36400 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_315
timestamp 1698431365
transform 1 0 36624 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_345
timestamp 1698431365
transform 1 0 39984 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_349
timestamp 1698431365
transform 1 0 40432 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_410
timestamp 1698431365
transform 1 0 47264 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_451
timestamp 1698431365
transform 1 0 51856 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_459
timestamp 1698431365
transform 1 0 52752 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_463
timestamp 1698431365
transform 1 0 53200 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698431365
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698431365
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698431365
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_107
timestamp 1698431365
transform 1 0 13328 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_115
timestamp 1698431365
transform 1 0 14224 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_145
timestamp 1698431365
transform 1 0 17584 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_149
timestamp 1698431365
transform 1 0 18032 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_153
timestamp 1698431365
transform 1 0 18480 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_161
timestamp 1698431365
transform 1 0 19376 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_169
timestamp 1698431365
transform 1 0 20272 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_173
timestamp 1698431365
transform 1 0 20720 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_177
timestamp 1698431365
transform 1 0 21168 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_185
timestamp 1698431365
transform 1 0 22064 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_193
timestamp 1698431365
transform 1 0 22960 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_201
timestamp 1698431365
transform 1 0 23856 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_205
timestamp 1698431365
transform 1 0 24304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_207
timestamp 1698431365
transform 1 0 24528 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_210
timestamp 1698431365
transform 1 0 24864 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_214
timestamp 1698431365
transform 1 0 25312 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_216
timestamp 1698431365
transform 1 0 25536 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_223
timestamp 1698431365
transform 1 0 26320 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_231
timestamp 1698431365
transform 1 0 27216 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_235
timestamp 1698431365
transform 1 0 27664 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_258
timestamp 1698431365
transform 1 0 30240 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_262
timestamp 1698431365
transform 1 0 30688 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_266
timestamp 1698431365
transform 1 0 31136 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_272
timestamp 1698431365
transform 1 0 31808 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_304
timestamp 1698431365
transform 1 0 35392 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_312
timestamp 1698431365
transform 1 0 36288 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_317
timestamp 1698431365
transform 1 0 36848 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_324
timestamp 1698431365
transform 1 0 37632 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_340
timestamp 1698431365
transform 1 0 39424 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_344
timestamp 1698431365
transform 1 0 39872 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_348
timestamp 1698431365
transform 1 0 40320 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_352
timestamp 1698431365
transform 1 0 40768 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_384
timestamp 1698431365
transform 1 0 44352 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_391
timestamp 1698431365
transform 1 0 45136 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_406
timestamp 1698431365
transform 1 0 46816 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_410
timestamp 1698431365
transform 1 0 47264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_414
timestamp 1698431365
transform 1 0 47712 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_424
timestamp 1698431365
transform 1 0 48832 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_428
timestamp 1698431365
transform 1 0 49280 0 1 4704
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_444
timestamp 1698431365
transform 1 0 51072 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_452
timestamp 1698431365
transform 1 0 51968 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_454
timestamp 1698431365
transform 1 0 52192 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_457
timestamp 1698431365
transform 1 0 52528 0 1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698431365
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698431365
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_72
timestamp 1698431365
transform 1 0 9408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_117
timestamp 1698431365
transform 1 0 14448 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_121
timestamp 1698431365
transform 1 0 14896 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_137
timestamp 1698431365
transform 1 0 16688 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_139
timestamp 1698431365
transform 1 0 16912 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_142
timestamp 1698431365
transform 1 0 17248 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_150
timestamp 1698431365
transform 1 0 18144 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_154
timestamp 1698431365
transform 1 0 18592 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_170
timestamp 1698431365
transform 1 0 20384 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_174
timestamp 1698431365
transform 1 0 20832 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_194
timestamp 1698431365
transform 1 0 23072 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_218
timestamp 1698431365
transform 1 0 25760 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_250
timestamp 1698431365
transform 1 0 29344 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_266
timestamp 1698431365
transform 1 0 31136 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_274
timestamp 1698431365
transform 1 0 32032 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_278
timestamp 1698431365
transform 1 0 32480 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_290
timestamp 1698431365
transform 1 0 33824 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_306
timestamp 1698431365
transform 1 0 35616 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_314
timestamp 1698431365
transform 1 0 36512 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_318
timestamp 1698431365
transform 1 0 36960 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_322
timestamp 1698431365
transform 1 0 37408 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_338
timestamp 1698431365
transform 1 0 39200 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_346
timestamp 1698431365
transform 1 0 40096 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_3_352
timestamp 1698431365
transform 1 0 40768 0 -1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_3_371
timestamp 1698431365
transform 1 0 42896 0 -1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_3_403
timestamp 1698431365
transform 1 0 46480 0 -1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_419
timestamp 1698431365
transform 1 0 48272 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_422
timestamp 1698431365
transform 1 0 48608 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_428
timestamp 1698431365
transform 1 0 49280 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698431365
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698431365
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_37
timestamp 1698431365
transform 1 0 5488 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_53
timestamp 1698431365
transform 1 0 7280 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_55
timestamp 1698431365
transform 1 0 7504 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_87
timestamp 1698431365
transform 1 0 11088 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_91
timestamp 1698431365
transform 1 0 11536 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_99
timestamp 1698431365
transform 1 0 12432 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_103
timestamp 1698431365
transform 1 0 12880 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_107
timestamp 1698431365
transform 1 0 13328 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_115
timestamp 1698431365
transform 1 0 14224 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_119
timestamp 1698431365
transform 1 0 14672 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_121
timestamp 1698431365
transform 1 0 14896 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_153
timestamp 1698431365
transform 1 0 18480 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_169
timestamp 1698431365
transform 1 0 20272 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_173
timestamp 1698431365
transform 1 0 20720 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_177
timestamp 1698431365
transform 1 0 21168 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_209
timestamp 1698431365
transform 1 0 24752 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_213
timestamp 1698431365
transform 1 0 25200 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_220
timestamp 1698431365
transform 1 0 25984 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_224
timestamp 1698431365
transform 1 0 26432 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_230
timestamp 1698431365
transform 1 0 27104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_237
timestamp 1698431365
transform 1 0 27888 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_247
timestamp 1698431365
transform 1 0 29008 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_254
timestamp 1698431365
transform 1 0 29792 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_317
timestamp 1698431365
transform 1 0 36848 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_332
timestamp 1698431365
transform 1 0 38528 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_336
timestamp 1698431365
transform 1 0 38976 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_4_340
timestamp 1698431365
transform 1 0 39424 0 1 6272
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_356
timestamp 1698431365
transform 1 0 41216 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_4_372
timestamp 1698431365
transform 1 0 43008 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_380
timestamp 1698431365
transform 1 0 43904 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_384
timestamp 1698431365
transform 1 0 44352 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_387
timestamp 1698431365
transform 1 0 44688 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_389
timestamp 1698431365
transform 1 0 44912 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_439
timestamp 1698431365
transform 1 0 50512 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_4_443
timestamp 1698431365
transform 1 0 50960 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_2
timestamp 1698431365
transform 1 0 1568 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_34
timestamp 1698431365
transform 1 0 5152 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_50
timestamp 1698431365
transform 1 0 6944 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_58
timestamp 1698431365
transform 1 0 7840 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_65
timestamp 1698431365
transform 1 0 8624 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_69
timestamp 1698431365
transform 1 0 9072 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_5_72
timestamp 1698431365
transform 1 0 9408 0 -1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_104
timestamp 1698431365
transform 1 0 12992 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_108
timestamp 1698431365
transform 1 0 13440 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_110
timestamp 1698431365
transform 1 0 13664 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_115
timestamp 1698431365
transform 1 0 14224 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_131
timestamp 1698431365
transform 1 0 16016 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_139
timestamp 1698431365
transform 1 0 16912 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_142
timestamp 1698431365
transform 1 0 17248 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_158
timestamp 1698431365
transform 1 0 19040 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_177
timestamp 1698431365
transform 1 0 21168 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_181
timestamp 1698431365
transform 1 0 21616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_189
timestamp 1698431365
transform 1 0 22512 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_193
timestamp 1698431365
transform 1 0 22960 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_201
timestamp 1698431365
transform 1 0 23856 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_209
timestamp 1698431365
transform 1 0 24752 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_212
timestamp 1698431365
transform 1 0 25088 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_228
timestamp 1698431365
transform 1 0 26880 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_236
timestamp 1698431365
transform 1 0 27776 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_244
timestamp 1698431365
transform 1 0 28672 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_252
timestamp 1698431365
transform 1 0 29568 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_260
timestamp 1698431365
transform 1 0 30464 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698431365
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_282
timestamp 1698431365
transform 1 0 32928 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_5_286
timestamp 1698431365
transform 1 0 33376 0 -1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_302
timestamp 1698431365
transform 1 0 35168 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_306
timestamp 1698431365
transform 1 0 35616 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_308
timestamp 1698431365
transform 1 0 35840 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_5_311
timestamp 1698431365
transform 1 0 36176 0 -1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_319
timestamp 1698431365
transform 1 0 37072 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_352
timestamp 1698431365
transform 1 0 40768 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_356
timestamp 1698431365
transform 1 0 41216 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_360
timestamp 1698431365
transform 1 0 41664 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_362
timestamp 1698431365
transform 1 0 41888 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_372
timestamp 1698431365
transform 1 0 43008 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_376
timestamp 1698431365
transform 1 0 43456 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_380
timestamp 1698431365
transform 1 0 43904 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_406
timestamp 1698431365
transform 1 0 46816 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_410
timestamp 1698431365
transform 1 0 47264 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_432
timestamp 1698431365
transform 1 0 49728 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698431365
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698431365
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_37
timestamp 1698431365
transform 1 0 5488 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_53
timestamp 1698431365
transform 1 0 7280 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_70
timestamp 1698431365
transform 1 0 9184 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_74
timestamp 1698431365
transform 1 0 9632 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_90
timestamp 1698431365
transform 1 0 11424 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_98
timestamp 1698431365
transform 1 0 12320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_102
timestamp 1698431365
transform 1 0 12768 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_104
timestamp 1698431365
transform 1 0 12992 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_107
timestamp 1698431365
transform 1 0 13328 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_111
timestamp 1698431365
transform 1 0 13776 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_127
timestamp 1698431365
transform 1 0 15568 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_135
timestamp 1698431365
transform 1 0 16464 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_139
timestamp 1698431365
transform 1 0 16912 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_142
timestamp 1698431365
transform 1 0 17248 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_158
timestamp 1698431365
transform 1 0 19040 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_177
timestamp 1698431365
transform 1 0 21168 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_181
timestamp 1698431365
transform 1 0 21616 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_221
timestamp 1698431365
transform 1 0 26096 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_225
timestamp 1698431365
transform 1 0 26544 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698431365
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_247
timestamp 1698431365
transform 1 0 29008 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_255
timestamp 1698431365
transform 1 0 29904 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_262
timestamp 1698431365
transform 1 0 30688 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_266
timestamp 1698431365
transform 1 0 31136 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_298
timestamp 1698431365
transform 1 0 34720 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_314
timestamp 1698431365
transform 1 0 36512 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_317
timestamp 1698431365
transform 1 0 36848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_325
timestamp 1698431365
transform 1 0 37744 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_332
timestamp 1698431365
transform 1 0 38528 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_348
timestamp 1698431365
transform 1 0 40320 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_365
timestamp 1698431365
transform 1 0 42224 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_6_369
timestamp 1698431365
transform 1 0 42672 0 1 7840
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_400
timestamp 1698431365
transform 1 0 46144 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_408
timestamp 1698431365
transform 1 0 47040 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_412
timestamp 1698431365
transform 1 0 47488 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_432
timestamp 1698431365
transform 1 0 49728 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_436
timestamp 1698431365
transform 1 0 50176 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_6_442
timestamp 1698431365
transform 1 0 50848 0 1 7840
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_450
timestamp 1698431365
transform 1 0 51744 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_454
timestamp 1698431365
transform 1 0 52192 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_6_463
timestamp 1698431365
transform 1 0 53200 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_2
timestamp 1698431365
transform 1 0 1568 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_18
timestamp 1698431365
transform 1 0 3360 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_55
timestamp 1698431365
transform 1 0 7504 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_59
timestamp 1698431365
transform 1 0 7952 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_67
timestamp 1698431365
transform 1 0 8848 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_69
timestamp 1698431365
transform 1 0 9072 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_72
timestamp 1698431365
transform 1 0 9408 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_74
timestamp 1698431365
transform 1 0 9632 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_137
timestamp 1698431365
transform 1 0 16688 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_139
timestamp 1698431365
transform 1 0 16912 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_7_171
timestamp 1698431365
transform 1 0 20496 0 -1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_203
timestamp 1698431365
transform 1 0 24080 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_207
timestamp 1698431365
transform 1 0 24528 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_209
timestamp 1698431365
transform 1 0 24752 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_212
timestamp 1698431365
transform 1 0 25088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_219
timestamp 1698431365
transform 1 0 25872 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_223
timestamp 1698431365
transform 1 0 26320 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_256
timestamp 1698431365
transform 1 0 30016 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_266
timestamp 1698431365
transform 1 0 31136 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_270
timestamp 1698431365
transform 1 0 31584 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_278
timestamp 1698431365
transform 1 0 32480 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_282
timestamp 1698431365
transform 1 0 32928 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_298
timestamp 1698431365
transform 1 0 34720 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_302
timestamp 1698431365
transform 1 0 35168 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_310
timestamp 1698431365
transform 1 0 36064 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_318
timestamp 1698431365
transform 1 0 36960 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_322
timestamp 1698431365
transform 1 0 37408 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_325
timestamp 1698431365
transform 1 0 37744 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_333
timestamp 1698431365
transform 1 0 38640 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_337
timestamp 1698431365
transform 1 0 39088 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_339
timestamp 1698431365
transform 1 0 39312 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_352
timestamp 1698431365
transform 1 0 40768 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_364
timestamp 1698431365
transform 1 0 42112 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_374
timestamp 1698431365
transform 1 0 43232 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_382
timestamp 1698431365
transform 1 0 44128 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_386
timestamp 1698431365
transform 1 0 44576 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_402
timestamp 1698431365
transform 1 0 46368 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_7_406
timestamp 1698431365
transform 1 0 46816 0 -1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_414
timestamp 1698431365
transform 1 0 47712 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_418
timestamp 1698431365
transform 1 0 48160 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_7_434
timestamp 1698431365
transform 1 0 49952 0 -1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_450
timestamp 1698431365
transform 1 0 51744 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_454
timestamp 1698431365
transform 1 0 52192 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_456
timestamp 1698431365
transform 1 0 52416 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698431365
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698431365
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_37
timestamp 1698431365
transform 1 0 5488 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_45
timestamp 1698431365
transform 1 0 6384 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_78
timestamp 1698431365
transform 1 0 10080 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_82
timestamp 1698431365
transform 1 0 10528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_90
timestamp 1698431365
transform 1 0 11424 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_96
timestamp 1698431365
transform 1 0 12096 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_104
timestamp 1698431365
transform 1 0 12992 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_107
timestamp 1698431365
transform 1 0 13328 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_123
timestamp 1698431365
transform 1 0 15120 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_127
timestamp 1698431365
transform 1 0 15568 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_133
timestamp 1698431365
transform 1 0 16240 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_139
timestamp 1698431365
transform 1 0 16912 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698431365
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_187
timestamp 1698431365
transform 1 0 22288 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_189
timestamp 1698431365
transform 1 0 22512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_8_195
timestamp 1698431365
transform 1 0 23184 0 1 9408
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_211
timestamp 1698431365
transform 1 0 24976 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_215
timestamp 1698431365
transform 1 0 25424 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_222
timestamp 1698431365
transform 1 0 26208 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_226
timestamp 1698431365
transform 1 0 26656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_230
timestamp 1698431365
transform 1 0 27104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_240
timestamp 1698431365
transform 1 0 28224 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_244
timestamp 1698431365
transform 1 0 28672 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_247
timestamp 1698431365
transform 1 0 29008 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_255
timestamp 1698431365
transform 1 0 29904 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_264
timestamp 1698431365
transform 1 0 30912 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_268
timestamp 1698431365
transform 1 0 31360 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_276
timestamp 1698431365
transform 1 0 32256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_278
timestamp 1698431365
transform 1 0 32480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_292
timestamp 1698431365
transform 1 0 34048 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_313
timestamp 1698431365
transform 1 0 36400 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_323
timestamp 1698431365
transform 1 0 37520 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_325
timestamp 1698431365
transform 1 0 37744 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_340
timestamp 1698431365
transform 1 0 39424 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_342
timestamp 1698431365
transform 1 0 39648 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_380
timestamp 1698431365
transform 1 0 43904 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_382
timestamp 1698431365
transform 1 0 44128 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_401
timestamp 1698431365
transform 1 0 46256 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_403
timestamp 1698431365
transform 1 0 46480 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_420
timestamp 1698431365
transform 1 0 48384 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_422
timestamp 1698431365
transform 1 0 48608 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_435
timestamp 1698431365
transform 1 0 50064 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_439
timestamp 1698431365
transform 1 0 50512 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_444
timestamp 1698431365
transform 1 0 51072 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_8_452
timestamp 1698431365
transform 1 0 51968 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_454
timestamp 1698431365
transform 1 0 52192 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_8_457
timestamp 1698431365
transform 1 0 52528 0 1 9408
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_31
timestamp 1698431365
transform 1 0 4816 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_35
timestamp 1698431365
transform 1 0 5264 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_67
timestamp 1698431365
transform 1 0 8848 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_69
timestamp 1698431365
transform 1 0 9072 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_72
timestamp 1698431365
transform 1 0 9408 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_80
timestamp 1698431365
transform 1 0 10304 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_104
timestamp 1698431365
transform 1 0 12992 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_108
timestamp 1698431365
transform 1 0 13440 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_142
timestamp 1698431365
transform 1 0 17248 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_158
timestamp 1698431365
transform 1 0 19040 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_166
timestamp 1698431365
transform 1 0 19936 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_170
timestamp 1698431365
transform 1 0 20384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_172
timestamp 1698431365
transform 1 0 20608 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_178
timestamp 1698431365
transform 1 0 21280 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_218
timestamp 1698431365
transform 1 0 25760 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_222
timestamp 1698431365
transform 1 0 26208 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_235
timestamp 1698431365
transform 1 0 27664 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_239
timestamp 1698431365
transform 1 0 28112 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_271
timestamp 1698431365
transform 1 0 31696 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_279
timestamp 1698431365
transform 1 0 32592 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_9_282
timestamp 1698431365
transform 1 0 32928 0 -1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_9_314
timestamp 1698431365
transform 1 0 36512 0 -1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_330
timestamp 1698431365
transform 1 0 38304 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_338
timestamp 1698431365
transform 1 0 39200 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_342
timestamp 1698431365
transform 1 0 39648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_346
timestamp 1698431365
transform 1 0 40096 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_352
timestamp 1698431365
transform 1 0 40768 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_361
timestamp 1698431365
transform 1 0 41776 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_365
timestamp 1698431365
transform 1 0 42224 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_372
timestamp 1698431365
transform 1 0 43008 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_376
timestamp 1698431365
transform 1 0 43456 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_380
timestamp 1698431365
transform 1 0 43904 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_398
timestamp 1698431365
transform 1 0 45920 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_400
timestamp 1698431365
transform 1 0 46144 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_9_411
timestamp 1698431365
transform 1 0 47376 0 -1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_419
timestamp 1698431365
transform 1 0 48272 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_422
timestamp 1698431365
transform 1 0 48608 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_2
timestamp 1698431365
transform 1 0 1568 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_18
timestamp 1698431365
transform 1 0 3360 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_26
timestamp 1698431365
transform 1 0 4256 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_30
timestamp 1698431365
transform 1 0 4704 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_48
timestamp 1698431365
transform 1 0 6720 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_52
timestamp 1698431365
transform 1 0 7168 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_56
timestamp 1698431365
transform 1 0 7616 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_73
timestamp 1698431365
transform 1 0 9520 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_81
timestamp 1698431365
transform 1 0 10416 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_91
timestamp 1698431365
transform 1 0 11536 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_99
timestamp 1698431365
transform 1 0 12432 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_103
timestamp 1698431365
transform 1 0 12880 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_107
timestamp 1698431365
transform 1 0 13328 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_111
timestamp 1698431365
transform 1 0 13776 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_132
timestamp 1698431365
transform 1 0 16128 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_167
timestamp 1698431365
transform 1 0 20048 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_177
timestamp 1698431365
transform 1 0 21168 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_207
timestamp 1698431365
transform 1 0 24528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_211
timestamp 1698431365
transform 1 0 24976 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_215
timestamp 1698431365
transform 1 0 25424 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_217
timestamp 1698431365
transform 1 0 25648 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_224
timestamp 1698431365
transform 1 0 26432 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_240
timestamp 1698431365
transform 1 0 28224 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_244
timestamp 1698431365
transform 1 0 28672 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_247
timestamp 1698431365
transform 1 0 29008 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_263
timestamp 1698431365
transform 1 0 30800 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_280
timestamp 1698431365
transform 1 0 32704 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_296
timestamp 1698431365
transform 1 0 34496 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_304
timestamp 1698431365
transform 1 0 35392 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_308
timestamp 1698431365
transform 1 0 35840 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_310
timestamp 1698431365
transform 1 0 36064 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_313
timestamp 1698431365
transform 1 0 36400 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_317
timestamp 1698431365
transform 1 0 36848 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_325
timestamp 1698431365
transform 1 0 37744 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_333
timestamp 1698431365
transform 1 0 38640 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_349
timestamp 1698431365
transform 1 0 40432 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_351
timestamp 1698431365
transform 1 0 40656 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_354
timestamp 1698431365
transform 1 0 40992 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_358
timestamp 1698431365
transform 1 0 41440 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_370
timestamp 1698431365
transform 1 0 42784 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_378
timestamp 1698431365
transform 1 0 43680 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_382
timestamp 1698431365
transform 1 0 44128 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_384
timestamp 1698431365
transform 1 0 44352 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_387
timestamp 1698431365
transform 1 0 44688 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_419
timestamp 1698431365
transform 1 0 48272 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_10_426
timestamp 1698431365
transform 1 0 49056 0 1 10976
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_10_436
timestamp 1698431365
transform 1 0 50176 0 1 10976
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_452
timestamp 1698431365
transform 1 0 51968 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_454
timestamp 1698431365
transform 1 0 52192 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_10_457
timestamp 1698431365
transform 1 0 52528 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_2
timestamp 1698431365
transform 1 0 1568 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_18
timestamp 1698431365
transform 1 0 3360 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_26
timestamp 1698431365
transform 1 0 4256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_30
timestamp 1698431365
transform 1 0 4704 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_33
timestamp 1698431365
transform 1 0 5040 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_49
timestamp 1698431365
transform 1 0 6832 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_67
timestamp 1698431365
transform 1 0 8848 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_69
timestamp 1698431365
transform 1 0 9072 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_72
timestamp 1698431365
transform 1 0 9408 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_74
timestamp 1698431365
transform 1 0 9632 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_85
timestamp 1698431365
transform 1 0 10864 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_93
timestamp 1698431365
transform 1 0 11760 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_105
timestamp 1698431365
transform 1 0 13104 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_109
timestamp 1698431365
transform 1 0 13552 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_122
timestamp 1698431365
transform 1 0 15008 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_138
timestamp 1698431365
transform 1 0 16800 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142
timestamp 1698431365
transform 1 0 17248 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_162
timestamp 1698431365
transform 1 0 19488 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_178
timestamp 1698431365
transform 1 0 21280 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_188
timestamp 1698431365
transform 1 0 22400 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_196
timestamp 1698431365
transform 1 0 23296 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_200
timestamp 1698431365
transform 1 0 23744 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_206
timestamp 1698431365
transform 1 0 24416 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_212
timestamp 1698431365
transform 1 0 25088 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_220
timestamp 1698431365
transform 1 0 25984 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_224
timestamp 1698431365
transform 1 0 26432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_238
timestamp 1698431365
transform 1 0 28000 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_242
timestamp 1698431365
transform 1 0 28448 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_244
timestamp 1698431365
transform 1 0 28672 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698431365
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_317
timestamp 1698431365
transform 1 0 36848 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_347
timestamp 1698431365
transform 1 0 40208 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_349
timestamp 1698431365
transform 1 0 40432 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_352
timestamp 1698431365
transform 1 0 40768 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_356
timestamp 1698431365
transform 1 0 41216 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_387
timestamp 1698431365
transform 1 0 44688 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_391
timestamp 1698431365
transform 1 0 45136 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_403
timestamp 1698431365
transform 1 0 46480 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_419
timestamp 1698431365
transform 1 0 48272 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_428
timestamp 1698431365
transform 1 0 49280 0 -1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_444
timestamp 1698431365
transform 1 0 51072 0 -1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_452
timestamp 1698431365
transform 1 0 51968 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_454
timestamp 1698431365
transform 1 0 52192 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_461
timestamp 1698431365
transform 1 0 52976 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_54
timestamp 1698431365
transform 1 0 7392 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_70
timestamp 1698431365
transform 1 0 9184 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_78
timestamp 1698431365
transform 1 0 10080 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_88
timestamp 1698431365
transform 1 0 11200 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_92
timestamp 1698431365
transform 1 0 11648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_96
timestamp 1698431365
transform 1 0 12096 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_104
timestamp 1698431365
transform 1 0 12992 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_107
timestamp 1698431365
transform 1 0 13328 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_121
timestamp 1698431365
transform 1 0 14896 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_131
timestamp 1698431365
transform 1 0 16016 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_147
timestamp 1698431365
transform 1 0 17808 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_158
timestamp 1698431365
transform 1 0 19040 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698431365
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698431365
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_189
timestamp 1698431365
transform 1 0 22512 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_197
timestamp 1698431365
transform 1 0 23408 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_201
timestamp 1698431365
transform 1 0 23856 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_207
timestamp 1698431365
transform 1 0 24528 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_211
timestamp 1698431365
transform 1 0 24976 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_213
timestamp 1698431365
transform 1 0 25200 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_247
timestamp 1698431365
transform 1 0 29008 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_279
timestamp 1698431365
transform 1 0 32592 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_295
timestamp 1698431365
transform 1 0 34384 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_303
timestamp 1698431365
transform 1 0 35280 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_314
timestamp 1698431365
transform 1 0 36512 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_317
timestamp 1698431365
transform 1 0 36848 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_325
timestamp 1698431365
transform 1 0 37744 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_336
timestamp 1698431365
transform 1 0 38976 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_352
timestamp 1698431365
transform 1 0 40768 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_360
timestamp 1698431365
transform 1 0 41664 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_367
timestamp 1698431365
transform 1 0 42448 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_375
timestamp 1698431365
transform 1 0 43344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_383
timestamp 1698431365
transform 1 0 44240 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_387
timestamp 1698431365
transform 1 0 44688 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_403
timestamp 1698431365
transform 1 0 46480 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_434
timestamp 1698431365
transform 1 0 49952 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_444
timestamp 1698431365
transform 1 0 51072 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_452
timestamp 1698431365
transform 1 0 51968 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_454
timestamp 1698431365
transform 1 0 52192 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_457
timestamp 1698431365
transform 1 0 52528 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_2
timestamp 1698431365
transform 1 0 1568 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_18
timestamp 1698431365
transform 1 0 3360 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_26
timestamp 1698431365
transform 1 0 4256 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_36
timestamp 1698431365
transform 1 0 5376 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_51
timestamp 1698431365
transform 1 0 7056 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_55
timestamp 1698431365
transform 1 0 7504 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_63
timestamp 1698431365
transform 1 0 8400 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_67
timestamp 1698431365
transform 1 0 8848 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_69
timestamp 1698431365
transform 1 0 9072 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_78
timestamp 1698431365
transform 1 0 10080 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_82
timestamp 1698431365
transform 1 0 10528 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_90
timestamp 1698431365
transform 1 0 11424 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_94
timestamp 1698431365
transform 1 0 11872 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_102
timestamp 1698431365
transform 1 0 12768 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_118
timestamp 1698431365
transform 1 0 14560 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_136
timestamp 1698431365
transform 1 0 16576 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698431365
transform 1 0 17248 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_146
timestamp 1698431365
transform 1 0 17696 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_166
timestamp 1698431365
transform 1 0 19936 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_170
timestamp 1698431365
transform 1 0 20384 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_207
timestamp 1698431365
transform 1 0 24528 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698431365
transform 1 0 24752 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698431365
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_216
timestamp 1698431365
transform 1 0 25536 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_224
timestamp 1698431365
transform 1 0 26432 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_226
timestamp 1698431365
transform 1 0 26656 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_258
timestamp 1698431365
transform 1 0 30240 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_266
timestamp 1698431365
transform 1 0 31136 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_270
timestamp 1698431365
transform 1 0 31584 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_282
timestamp 1698431365
transform 1 0 32928 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_286
timestamp 1698431365
transform 1 0 33376 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_293
timestamp 1698431365
transform 1 0 34160 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_313
timestamp 1698431365
transform 1 0 36400 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_329
timestamp 1698431365
transform 1 0 38192 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_337
timestamp 1698431365
transform 1 0 39088 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_347
timestamp 1698431365
transform 1 0 40208 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_349
timestamp 1698431365
transform 1 0 40432 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_352
timestamp 1698431365
transform 1 0 40768 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_416
timestamp 1698431365
transform 1 0 47936 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_422
timestamp 1698431365
transform 1 0 48608 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_430
timestamp 1698431365
transform 1 0 49504 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698431365
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698431365
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_37
timestamp 1698431365
transform 1 0 5488 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_45
timestamp 1698431365
transform 1 0 6384 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_57
timestamp 1698431365
transform 1 0 7728 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_61
timestamp 1698431365
transform 1 0 8176 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_63
timestamp 1698431365
transform 1 0 8400 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_66
timestamp 1698431365
transform 1 0 8736 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_74
timestamp 1698431365
transform 1 0 9632 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_84
timestamp 1698431365
transform 1 0 10752 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_97
timestamp 1698431365
transform 1 0 12208 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_107
timestamp 1698431365
transform 1 0 13328 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_147
timestamp 1698431365
transform 1 0 17808 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_151
timestamp 1698431365
transform 1 0 18256 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_153
timestamp 1698431365
transform 1 0 18480 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_160
timestamp 1698431365
transform 1 0 19264 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_168
timestamp 1698431365
transform 1 0 20160 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698431365
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698431365
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698431365
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698431365
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_189
timestamp 1698431365
transform 1 0 22512 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_199
timestamp 1698431365
transform 1 0 23632 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_207
timestamp 1698431365
transform 1 0 24528 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_223
timestamp 1698431365
transform 1 0 26320 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_227
timestamp 1698431365
transform 1 0 26768 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698431365
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_247
timestamp 1698431365
transform 1 0 29008 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_263
timestamp 1698431365
transform 1 0 30800 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_271
timestamp 1698431365
transform 1 0 31696 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_286
timestamp 1698431365
transform 1 0 33376 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_294
timestamp 1698431365
transform 1 0 34272 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_296
timestamp 1698431365
transform 1 0 34496 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_299
timestamp 1698431365
transform 1 0 34832 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_301
timestamp 1698431365
transform 1 0 35056 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_310
timestamp 1698431365
transform 1 0 36064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_314
timestamp 1698431365
transform 1 0 36512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_317
timestamp 1698431365
transform 1 0 36848 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_325
timestamp 1698431365
transform 1 0 37744 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_339
timestamp 1698431365
transform 1 0 39312 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_347
timestamp 1698431365
transform 1 0 40208 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_358
timestamp 1698431365
transform 1 0 41440 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_360
timestamp 1698431365
transform 1 0 41664 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_367
timestamp 1698431365
transform 1 0 42448 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_377
timestamp 1698431365
transform 1 0 43568 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_387
timestamp 1698431365
transform 1 0 44688 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_395
timestamp 1698431365
transform 1 0 45584 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_397
timestamp 1698431365
transform 1 0 45808 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_404
timestamp 1698431365
transform 1 0 46592 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_408
timestamp 1698431365
transform 1 0 47040 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_416
timestamp 1698431365
transform 1 0 47936 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_428
timestamp 1698431365
transform 1 0 49280 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_444
timestamp 1698431365
transform 1 0 51072 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_452
timestamp 1698431365
transform 1 0 51968 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_2
timestamp 1698431365
transform 1 0 1568 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_6
timestamp 1698431365
transform 1 0 2016 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_13
timestamp 1698431365
transform 1 0 2800 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_21
timestamp 1698431365
transform 1 0 3696 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_25
timestamp 1698431365
transform 1 0 4144 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_27
timestamp 1698431365
transform 1 0 4368 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_34
timestamp 1698431365
transform 1 0 5152 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_42
timestamp 1698431365
transform 1 0 6048 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_46
timestamp 1698431365
transform 1 0 6496 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_48
timestamp 1698431365
transform 1 0 6720 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_69
timestamp 1698431365
transform 1 0 9072 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_72
timestamp 1698431365
transform 1 0 9408 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_76
timestamp 1698431365
transform 1 0 9856 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698431365
transform 1 0 11648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698431365
transform 1 0 11872 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_133
timestamp 1698431365
transform 1 0 16240 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698431365
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698431365
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_142
timestamp 1698431365
transform 1 0 17248 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_150
timestamp 1698431365
transform 1 0 18144 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_161
timestamp 1698431365
transform 1 0 19376 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_165
timestamp 1698431365
transform 1 0 19824 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_169
timestamp 1698431365
transform 1 0 20272 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_175
timestamp 1698431365
transform 1 0 20944 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_183
timestamp 1698431365
transform 1 0 21840 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698431365
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_216
timestamp 1698431365
transform 1 0 25536 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_257
timestamp 1698431365
transform 1 0 30128 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_259
timestamp 1698431365
transform 1 0 30352 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_274
timestamp 1698431365
transform 1 0 32032 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698431365
transform 1 0 32480 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_282
timestamp 1698431365
transform 1 0 32928 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_290
timestamp 1698431365
transform 1 0 33824 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_346
timestamp 1698431365
transform 1 0 40096 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_352
timestamp 1698431365
transform 1 0 40768 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_360
timestamp 1698431365
transform 1 0 41664 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_371
timestamp 1698431365
transform 1 0 42896 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_389
timestamp 1698431365
transform 1 0 44912 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_397
timestamp 1698431365
transform 1 0 45808 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_401
timestamp 1698431365
transform 1 0 46256 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_410
timestamp 1698431365
transform 1 0 47264 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_414
timestamp 1698431365
transform 1 0 47712 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_418
timestamp 1698431365
transform 1 0 48160 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_427
timestamp 1698431365
transform 1 0 49168 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_442
timestamp 1698431365
transform 1 0 50848 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_458
timestamp 1698431365
transform 1 0 52640 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_462
timestamp 1698431365
transform 1 0 53088 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_31
timestamp 1698431365
transform 1 0 4816 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_37
timestamp 1698431365
transform 1 0 5488 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_39
timestamp 1698431365
transform 1 0 5712 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_48
timestamp 1698431365
transform 1 0 6720 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_60
timestamp 1698431365
transform 1 0 8064 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_68
timestamp 1698431365
transform 1 0 8960 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_72
timestamp 1698431365
transform 1 0 9408 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_74
timestamp 1698431365
transform 1 0 9632 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_85
timestamp 1698431365
transform 1 0 10864 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_89
timestamp 1698431365
transform 1 0 11312 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_95
timestamp 1698431365
transform 1 0 11984 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_99
timestamp 1698431365
transform 1 0 12432 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_103
timestamp 1698431365
transform 1 0 12880 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698431365
transform 1 0 13328 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_129
timestamp 1698431365
transform 1 0 15792 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_141
timestamp 1698431365
transform 1 0 17136 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_148
timestamp 1698431365
transform 1 0 17920 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_152
timestamp 1698431365
transform 1 0 18368 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_168
timestamp 1698431365
transform 1 0 20160 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698431365
transform 1 0 20608 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698431365
transform 1 0 20832 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_177
timestamp 1698431365
transform 1 0 21168 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_183
timestamp 1698431365
transform 1 0 21840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_187
timestamp 1698431365
transform 1 0 22288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_218
timestamp 1698431365
transform 1 0 25760 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_222
timestamp 1698431365
transform 1 0 26208 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_238
timestamp 1698431365
transform 1 0 28000 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698431365
transform 1 0 28448 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698431365
transform 1 0 28672 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_247
timestamp 1698431365
transform 1 0 29008 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_279
timestamp 1698431365
transform 1 0 32592 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_284
timestamp 1698431365
transform 1 0 33152 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_292
timestamp 1698431365
transform 1 0 34048 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_296
timestamp 1698431365
transform 1 0 34496 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_298
timestamp 1698431365
transform 1 0 34720 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_301
timestamp 1698431365
transform 1 0 35056 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_309
timestamp 1698431365
transform 1 0 35952 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_313
timestamp 1698431365
transform 1 0 36400 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_317
timestamp 1698431365
transform 1 0 36848 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_321
timestamp 1698431365
transform 1 0 37296 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_373
timestamp 1698431365
transform 1 0 43120 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_381
timestamp 1698431365
transform 1 0 44016 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_416
timestamp 1698431365
transform 1 0 47936 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_426
timestamp 1698431365
transform 1 0 49056 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_438
timestamp 1698431365
transform 1 0 50400 0 1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_454
timestamp 1698431365
transform 1 0 52192 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_457
timestamp 1698431365
transform 1 0 52528 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_2
timestamp 1698431365
transform 1 0 1568 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_18
timestamp 1698431365
transform 1 0 3360 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_26
timestamp 1698431365
transform 1 0 4256 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_33
timestamp 1698431365
transform 1 0 5040 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_65
timestamp 1698431365
transform 1 0 8624 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_69
timestamp 1698431365
transform 1 0 9072 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_111
timestamp 1698431365
transform 1 0 13776 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_115
timestamp 1698431365
transform 1 0 14224 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_126
timestamp 1698431365
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698431365
transform 1 0 16800 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_181
timestamp 1698431365
transform 1 0 21616 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_183
timestamp 1698431365
transform 1 0 21840 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698431365
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_216
timestamp 1698431365
transform 1 0 25536 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_282
timestamp 1698431365
transform 1 0 32928 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_284
timestamp 1698431365
transform 1 0 33152 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_333
timestamp 1698431365
transform 1 0 38640 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_337
timestamp 1698431365
transform 1 0 39088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_345
timestamp 1698431365
transform 1 0 39984 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_349
timestamp 1698431365
transform 1 0 40432 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_352
timestamp 1698431365
transform 1 0 40768 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_372
timestamp 1698431365
transform 1 0 43008 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_404
timestamp 1698431365
transform 1 0 46592 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_427
timestamp 1698431365
transform 1 0 49168 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_2
timestamp 1698431365
transform 1 0 1568 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_18
timestamp 1698431365
transform 1 0 3360 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_26
timestamp 1698431365
transform 1 0 4256 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_30
timestamp 1698431365
transform 1 0 4704 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_33
timestamp 1698431365
transform 1 0 5040 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_37
timestamp 1698431365
transform 1 0 5488 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_39
timestamp 1698431365
transform 1 0 5712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_50
timestamp 1698431365
transform 1 0 6944 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_54
timestamp 1698431365
transform 1 0 7392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_61
timestamp 1698431365
transform 1 0 8176 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_93
timestamp 1698431365
transform 1 0 11760 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698431365
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698431365
transform 1 0 13328 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698431365
transform 1 0 14224 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_119
timestamp 1698431365
transform 1 0 14672 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_121
timestamp 1698431365
transform 1 0 14896 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1698431365
transform 1 0 15456 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_130
timestamp 1698431365
transform 1 0 15904 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_162
timestamp 1698431365
transform 1 0 19488 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_170
timestamp 1698431365
transform 1 0 20384 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698431365
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_185
timestamp 1698431365
transform 1 0 22064 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_193
timestamp 1698431365
transform 1 0 22960 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_195
timestamp 1698431365
transform 1 0 23184 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_201
timestamp 1698431365
transform 1 0 23856 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_233
timestamp 1698431365
transform 1 0 27440 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698431365
transform 1 0 28336 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_247
timestamp 1698431365
transform 1 0 29008 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_251
timestamp 1698431365
transform 1 0 29456 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_289
timestamp 1698431365
transform 1 0 33712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_294
timestamp 1698431365
transform 1 0 34272 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_310
timestamp 1698431365
transform 1 0 36064 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_317
timestamp 1698431365
transform 1 0 36848 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_376
timestamp 1698431365
transform 1 0 43456 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_384
timestamp 1698431365
transform 1 0 44352 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_387
timestamp 1698431365
transform 1 0 44688 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_403
timestamp 1698431365
transform 1 0 46480 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_411
timestamp 1698431365
transform 1 0 47376 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_422
timestamp 1698431365
transform 1 0 48608 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_426
timestamp 1698431365
transform 1 0 49056 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_435
timestamp 1698431365
transform 1 0 50064 0 1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_451
timestamp 1698431365
transform 1 0 51856 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_457
timestamp 1698431365
transform 1 0 52528 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_48
timestamp 1698431365
transform 1 0 6720 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_52
timestamp 1698431365
transform 1 0 7168 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_54
timestamp 1698431365
transform 1 0 7392 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_57
timestamp 1698431365
transform 1 0 7728 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_65
timestamp 1698431365
transform 1 0 8624 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_69
timestamp 1698431365
transform 1 0 9072 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698431365
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698431365
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_121
timestamp 1698431365
transform 1 0 14896 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_125
timestamp 1698431365
transform 1 0 15344 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_133
timestamp 1698431365
transform 1 0 16240 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_137
timestamp 1698431365
transform 1 0 16688 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698431365
transform 1 0 16912 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_142
timestamp 1698431365
transform 1 0 17248 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_150
timestamp 1698431365
transform 1 0 18144 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_155
timestamp 1698431365
transform 1 0 18704 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_163
timestamp 1698431365
transform 1 0 19600 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_193
timestamp 1698431365
transform 1 0 22960 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_197
timestamp 1698431365
transform 1 0 23408 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_205
timestamp 1698431365
transform 1 0 24304 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698431365
transform 1 0 24752 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_217
timestamp 1698431365
transform 1 0 25648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_252
timestamp 1698431365
transform 1 0 29568 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_268
timestamp 1698431365
transform 1 0 31360 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_276
timestamp 1698431365
transform 1 0 32256 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_282
timestamp 1698431365
transform 1 0 32928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_286
timestamp 1698431365
transform 1 0 33376 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_333
timestamp 1698431365
transform 1 0 38640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_337
timestamp 1698431365
transform 1 0 39088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_345
timestamp 1698431365
transform 1 0 39984 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_349
timestamp 1698431365
transform 1 0 40432 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_352
timestamp 1698431365
transform 1 0 40768 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_360
timestamp 1698431365
transform 1 0 41664 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_392
timestamp 1698431365
transform 1 0 45248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_407
timestamp 1698431365
transform 1 0 46928 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_411
timestamp 1698431365
transform 1 0 47376 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_419
timestamp 1698431365
transform 1 0 48272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_422
timestamp 1698431365
transform 1 0 48608 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_430
timestamp 1698431365
transform 1 0 49504 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_440
timestamp 1698431365
transform 1 0 50624 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_447
timestamp 1698431365
transform 1 0 51408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_2
timestamp 1698431365
transform 1 0 1568 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_18
timestamp 1698431365
transform 1 0 3360 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_26
timestamp 1698431365
transform 1 0 4256 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_61
timestamp 1698431365
transform 1 0 8176 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_63
timestamp 1698431365
transform 1 0 8400 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_66
timestamp 1698431365
transform 1 0 8736 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_70
timestamp 1698431365
transform 1 0 9184 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_74
timestamp 1698431365
transform 1 0 9632 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_76
timestamp 1698431365
transform 1 0 9856 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_83
timestamp 1698431365
transform 1 0 10640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_93
timestamp 1698431365
transform 1 0 11760 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_97
timestamp 1698431365
transform 1 0 12208 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698431365
transform 1 0 13328 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698431365
transform 1 0 15120 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_156
timestamp 1698431365
transform 1 0 18816 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_172
timestamp 1698431365
transform 1 0 20608 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698431365
transform 1 0 20832 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_177
timestamp 1698431365
transform 1 0 21168 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_185
timestamp 1698431365
transform 1 0 22064 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_223
timestamp 1698431365
transform 1 0 26320 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_239
timestamp 1698431365
transform 1 0 28112 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698431365
transform 1 0 28560 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_247
timestamp 1698431365
transform 1 0 29008 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_255
timestamp 1698431365
transform 1 0 29904 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_273
timestamp 1698431365
transform 1 0 31920 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_287
timestamp 1698431365
transform 1 0 33488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698431365
transform 1 0 35840 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698431365
transform 1 0 36288 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698431365
transform 1 0 36512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_317
timestamp 1698431365
transform 1 0 36848 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_325
timestamp 1698431365
transform 1 0 37744 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_329
timestamp 1698431365
transform 1 0 38192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_348
timestamp 1698431365
transform 1 0 40320 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_356
timestamp 1698431365
transform 1 0 41216 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_362
timestamp 1698431365
transform 1 0 41888 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_366
timestamp 1698431365
transform 1 0 42336 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_382
timestamp 1698431365
transform 1 0 44128 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_384
timestamp 1698431365
transform 1 0 44352 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_387
timestamp 1698431365
transform 1 0 44688 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_395
timestamp 1698431365
transform 1 0 45584 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_397
timestamp 1698431365
transform 1 0 45808 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_406
timestamp 1698431365
transform 1 0 46816 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_439
timestamp 1698431365
transform 1 0 50512 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_446
timestamp 1698431365
transform 1 0 51296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_454
timestamp 1698431365
transform 1 0 52192 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_457
timestamp 1698431365
transform 1 0 52528 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_2
timestamp 1698431365
transform 1 0 1568 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_34
timestamp 1698431365
transform 1 0 5152 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_38
timestamp 1698431365
transform 1 0 5600 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_40
timestamp 1698431365
transform 1 0 5824 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_56
timestamp 1698431365
transform 1 0 7616 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_72
timestamp 1698431365
transform 1 0 9408 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_80
timestamp 1698431365
transform 1 0 10304 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_112
timestamp 1698431365
transform 1 0 13888 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_134
timestamp 1698431365
transform 1 0 16352 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698431365
transform 1 0 16800 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_142
timestamp 1698431365
transform 1 0 17248 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_150
timestamp 1698431365
transform 1 0 18144 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_158
timestamp 1698431365
transform 1 0 19040 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_190
timestamp 1698431365
transform 1 0 22624 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_206
timestamp 1698431365
transform 1 0 24416 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_220
timestamp 1698431365
transform 1 0 25984 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_228
timestamp 1698431365
transform 1 0 26880 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_232
timestamp 1698431365
transform 1 0 27328 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_234
timestamp 1698431365
transform 1 0 27552 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_247
timestamp 1698431365
transform 1 0 29008 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_251
timestamp 1698431365
transform 1 0 29456 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_255
timestamp 1698431365
transform 1 0 29904 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_258
timestamp 1698431365
transform 1 0 30240 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_260
timestamp 1698431365
transform 1 0 30464 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_263
timestamp 1698431365
transform 1 0 30800 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_279
timestamp 1698431365
transform 1 0 32592 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698431365
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_314
timestamp 1698431365
transform 1 0 36512 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_330
timestamp 1698431365
transform 1 0 38304 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_338
timestamp 1698431365
transform 1 0 39200 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_360
timestamp 1698431365
transform 1 0 41664 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_362
timestamp 1698431365
transform 1 0 41888 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_408
timestamp 1698431365
transform 1 0 47040 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_416
timestamp 1698431365
transform 1 0 47936 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_422
timestamp 1698431365
transform 1 0 48608 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_434
timestamp 1698431365
transform 1 0 49952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698431365
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698431365
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_37
timestamp 1698431365
transform 1 0 5488 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_53
timestamp 1698431365
transform 1 0 7280 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_60
timestamp 1698431365
transform 1 0 8064 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_86
timestamp 1698431365
transform 1 0 10976 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_102
timestamp 1698431365
transform 1 0 12768 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698431365
transform 1 0 12992 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698431365
transform 1 0 13328 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_109
timestamp 1698431365
transform 1 0 13552 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_122
timestamp 1698431365
transform 1 0 15008 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_161
timestamp 1698431365
transform 1 0 19376 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_168
timestamp 1698431365
transform 1 0 20160 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_172
timestamp 1698431365
transform 1 0 20608 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698431365
transform 1 0 20832 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_177
timestamp 1698431365
transform 1 0 21168 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_181
timestamp 1698431365
transform 1 0 21616 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_188
timestamp 1698431365
transform 1 0 22400 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_220
timestamp 1698431365
transform 1 0 25984 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698431365
transform 1 0 28672 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_252
timestamp 1698431365
transform 1 0 29568 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_256
timestamp 1698431365
transform 1 0 30016 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_292
timestamp 1698431365
transform 1 0 34048 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_308
timestamp 1698431365
transform 1 0 35840 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_312
timestamp 1698431365
transform 1 0 36288 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_314
timestamp 1698431365
transform 1 0 36512 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_317
timestamp 1698431365
transform 1 0 36848 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_333
timestamp 1698431365
transform 1 0 38640 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_337
timestamp 1698431365
transform 1 0 39088 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_384
timestamp 1698431365
transform 1 0 44352 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_391
timestamp 1698431365
transform 1 0 45136 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_395
timestamp 1698431365
transform 1 0 45584 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_405
timestamp 1698431365
transform 1 0 46704 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_409
timestamp 1698431365
transform 1 0 47152 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_413
timestamp 1698431365
transform 1 0 47600 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_429
timestamp 1698431365
transform 1 0 49392 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_433
timestamp 1698431365
transform 1 0 49840 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_436
timestamp 1698431365
transform 1 0 50176 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_452
timestamp 1698431365
transform 1 0 51968 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_454
timestamp 1698431365
transform 1 0 52192 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_457
timestamp 1698431365
transform 1 0 52528 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_31
timestamp 1698431365
transform 1 0 4816 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_37
timestamp 1698431365
transform 1 0 5488 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_41
timestamp 1698431365
transform 1 0 5936 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_57
timestamp 1698431365
transform 1 0 7728 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_63
timestamp 1698431365
transform 1 0 8400 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_67
timestamp 1698431365
transform 1 0 8848 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_69
timestamp 1698431365
transform 1 0 9072 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_72
timestamp 1698431365
transform 1 0 9408 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698431365
transform 1 0 13776 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_115
timestamp 1698431365
transform 1 0 14224 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_119
timestamp 1698431365
transform 1 0 14672 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_121
timestamp 1698431365
transform 1 0 14896 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_124
timestamp 1698431365
transform 1 0 15232 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_128
timestamp 1698431365
transform 1 0 15680 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_136
timestamp 1698431365
transform 1 0 16576 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_142
timestamp 1698431365
transform 1 0 17248 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_174
timestamp 1698431365
transform 1 0 20832 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_178
timestamp 1698431365
transform 1 0 21280 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_185
timestamp 1698431365
transform 1 0 22064 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_203
timestamp 1698431365
transform 1 0 24080 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698431365
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698431365
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_212
timestamp 1698431365
transform 1 0 25088 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698431365
transform 1 0 32256 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_282
timestamp 1698431365
transform 1 0 32928 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_292
timestamp 1698431365
transform 1 0 34048 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_296
timestamp 1698431365
transform 1 0 34496 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_300
timestamp 1698431365
transform 1 0 34944 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_330
timestamp 1698431365
transform 1 0 38304 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_334
timestamp 1698431365
transform 1 0 38752 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_338
timestamp 1698431365
transform 1 0 39200 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_349
timestamp 1698431365
transform 1 0 40432 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_358
timestamp 1698431365
transform 1 0 41440 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_362
timestamp 1698431365
transform 1 0 41888 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_366
timestamp 1698431365
transform 1 0 42336 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_383
timestamp 1698431365
transform 1 0 44240 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_387
timestamp 1698431365
transform 1 0 44688 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_391
timestamp 1698431365
transform 1 0 45136 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_395
timestamp 1698431365
transform 1 0 45584 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_418
timestamp 1698431365
transform 1 0 48160 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_432
timestamp 1698431365
transform 1 0 49728 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_436
timestamp 1698431365
transform 1 0 50176 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_440
timestamp 1698431365
transform 1 0 50624 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_456
timestamp 1698431365
transform 1 0 52416 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_460
timestamp 1698431365
transform 1 0 52864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_462
timestamp 1698431365
transform 1 0 53088 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_2
timestamp 1698431365
transform 1 0 1568 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_18
timestamp 1698431365
transform 1 0 3360 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_26
timestamp 1698431365
transform 1 0 4256 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_28
timestamp 1698431365
transform 1 0 4480 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_45
timestamp 1698431365
transform 1 0 6384 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_49
timestamp 1698431365
transform 1 0 6832 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_65
timestamp 1698431365
transform 1 0 8624 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_69
timestamp 1698431365
transform 1 0 9072 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_72
timestamp 1698431365
transform 1 0 9408 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_104
timestamp 1698431365
transform 1 0 12992 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_107
timestamp 1698431365
transform 1 0 13328 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_171
timestamp 1698431365
transform 1 0 20496 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_177
timestamp 1698431365
transform 1 0 21168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_184
timestamp 1698431365
transform 1 0 21952 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_200
timestamp 1698431365
transform 1 0 23744 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_226
timestamp 1698431365
transform 1 0 26656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_230
timestamp 1698431365
transform 1 0 27104 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_242
timestamp 1698431365
transform 1 0 28448 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698431365
transform 1 0 28672 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_247
timestamp 1698431365
transform 1 0 29008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_253
timestamp 1698431365
transform 1 0 29680 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_285
timestamp 1698431365
transform 1 0 33264 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_289
timestamp 1698431365
transform 1 0 33712 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_298
timestamp 1698431365
transform 1 0 34720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_310
timestamp 1698431365
transform 1 0 36064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698431365
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_322
timestamp 1698431365
transform 1 0 37408 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_326
timestamp 1698431365
transform 1 0 37856 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_363
timestamp 1698431365
transform 1 0 42000 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_381
timestamp 1698431365
transform 1 0 44016 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_387
timestamp 1698431365
transform 1 0 44688 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_421
timestamp 1698431365
transform 1 0 48496 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_427
timestamp 1698431365
transform 1 0 49168 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_447
timestamp 1698431365
transform 1 0 51408 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_457
timestamp 1698431365
transform 1 0 52528 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_2
timestamp 1698431365
transform 1 0 1568 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_6
timestamp 1698431365
transform 1 0 2016 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_8
timestamp 1698431365
transform 1 0 2240 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_15
timestamp 1698431365
transform 1 0 3024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_19
timestamp 1698431365
transform 1 0 3472 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_46
timestamp 1698431365
transform 1 0 6496 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_50
timestamp 1698431365
transform 1 0 6944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_60
timestamp 1698431365
transform 1 0 8064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_87
timestamp 1698431365
transform 1 0 11088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_91
timestamp 1698431365
transform 1 0 11536 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_95
timestamp 1698431365
transform 1 0 11984 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_97
timestamp 1698431365
transform 1 0 12208 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_129
timestamp 1698431365
transform 1 0 15792 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_137
timestamp 1698431365
transform 1 0 16688 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698431365
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_142
timestamp 1698431365
transform 1 0 17248 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_158
timestamp 1698431365
transform 1 0 19040 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_161
timestamp 1698431365
transform 1 0 19376 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_169
timestamp 1698431365
transform 1 0 20272 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_173
timestamp 1698431365
transform 1 0 20720 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_177
timestamp 1698431365
transform 1 0 21168 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_185
timestamp 1698431365
transform 1 0 22064 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_195
timestamp 1698431365
transform 1 0 23184 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_203
timestamp 1698431365
transform 1 0 24080 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_207
timestamp 1698431365
transform 1 0 24528 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698431365
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_212
timestamp 1698431365
transform 1 0 25088 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_220
timestamp 1698431365
transform 1 0 25984 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_252
timestamp 1698431365
transform 1 0 29568 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_260
timestamp 1698431365
transform 1 0 30464 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_274
timestamp 1698431365
transform 1 0 32032 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_278
timestamp 1698431365
transform 1 0 32480 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_282
timestamp 1698431365
transform 1 0 32928 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_300
timestamp 1698431365
transform 1 0 34944 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_304
timestamp 1698431365
transform 1 0 35392 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_312
timestamp 1698431365
transform 1 0 36288 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_314
timestamp 1698431365
transform 1 0 36512 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_317
timestamp 1698431365
transform 1 0 36848 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_321
timestamp 1698431365
transform 1 0 37296 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_348
timestamp 1698431365
transform 1 0 40320 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_352
timestamp 1698431365
transform 1 0 40768 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_388
timestamp 1698431365
transform 1 0 44800 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_427
timestamp 1698431365
transform 1 0 49168 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_31
timestamp 1698431365
transform 1 0 4816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_51
timestamp 1698431365
transform 1 0 7056 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_53
timestamp 1698431365
transform 1 0 7280 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_63
timestamp 1698431365
transform 1 0 8400 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_73
timestamp 1698431365
transform 1 0 9520 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698431365
transform 1 0 13328 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_123
timestamp 1698431365
transform 1 0 15120 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_130
timestamp 1698431365
transform 1 0 15904 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_138
timestamp 1698431365
transform 1 0 16800 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_142
timestamp 1698431365
transform 1 0 17248 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698431365
transform 1 0 21168 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_179
timestamp 1698431365
transform 1 0 21392 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_211
timestamp 1698431365
transform 1 0 24976 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698431365
transform 1 0 26320 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_227
timestamp 1698431365
transform 1 0 26768 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_240
timestamp 1698431365
transform 1 0 28224 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698431365
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_247
timestamp 1698431365
transform 1 0 29008 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_269
timestamp 1698431365
transform 1 0 31472 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_277
timestamp 1698431365
transform 1 0 32368 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_283
timestamp 1698431365
transform 1 0 33040 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_287
timestamp 1698431365
transform 1 0 33488 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_289
timestamp 1698431365
transform 1 0 33712 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_302
timestamp 1698431365
transform 1 0 35168 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_310
timestamp 1698431365
transform 1 0 36064 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_314
timestamp 1698431365
transform 1 0 36512 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698431365
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_328
timestamp 1698431365
transform 1 0 38080 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_332
timestamp 1698431365
transform 1 0 38528 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_338
timestamp 1698431365
transform 1 0 39200 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_346
timestamp 1698431365
transform 1 0 40096 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_348
timestamp 1698431365
transform 1 0 40320 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_379
timestamp 1698431365
transform 1 0 43792 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_383
timestamp 1698431365
transform 1 0 44240 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_387
timestamp 1698431365
transform 1 0 44688 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_391
timestamp 1698431365
transform 1 0 45136 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_415
timestamp 1698431365
transform 1 0 47824 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_447
timestamp 1698431365
transform 1 0 51408 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_457
timestamp 1698431365
transform 1 0 52528 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_2
timestamp 1698431365
transform 1 0 1568 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_18
timestamp 1698431365
transform 1 0 3360 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_26
timestamp 1698431365
transform 1 0 4256 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_38
timestamp 1698431365
transform 1 0 5600 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_72
timestamp 1698431365
transform 1 0 9408 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_76
timestamp 1698431365
transform 1 0 9856 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_119
timestamp 1698431365
transform 1 0 14672 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_127
timestamp 1698431365
transform 1 0 15568 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698431365
transform 1 0 17248 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_159
timestamp 1698431365
transform 1 0 19152 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_174
timestamp 1698431365
transform 1 0 20832 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_178
timestamp 1698431365
transform 1 0 21280 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_182
timestamp 1698431365
transform 1 0 21728 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_195
timestamp 1698431365
transform 1 0 23184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698431365
transform 1 0 23632 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_207
timestamp 1698431365
transform 1 0 24528 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698431365
transform 1 0 25088 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_216
timestamp 1698431365
transform 1 0 25536 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_225
timestamp 1698431365
transform 1 0 26544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_229
timestamp 1698431365
transform 1 0 26992 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_237
timestamp 1698431365
transform 1 0 27888 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_241
timestamp 1698431365
transform 1 0 28336 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_243
timestamp 1698431365
transform 1 0 28560 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_249
timestamp 1698431365
transform 1 0 29232 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698431365
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_282
timestamp 1698431365
transform 1 0 32928 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_317
timestamp 1698431365
transform 1 0 36848 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_321
timestamp 1698431365
transform 1 0 37296 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_352
timestamp 1698431365
transform 1 0 40768 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_360
timestamp 1698431365
transform 1 0 41664 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_364
timestamp 1698431365
transform 1 0 42112 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_367
timestamp 1698431365
transform 1 0 42448 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_378
timestamp 1698431365
transform 1 0 43680 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_382
timestamp 1698431365
transform 1 0 44128 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_390
timestamp 1698431365
transform 1 0 45024 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_394
timestamp 1698431365
transform 1 0 45472 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_404
timestamp 1698431365
transform 1 0 46592 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_422
timestamp 1698431365
transform 1 0 48608 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_438
timestamp 1698431365
transform 1 0 50400 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_442
timestamp 1698431365
transform 1 0 50848 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_458
timestamp 1698431365
transform 1 0 52640 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_462
timestamp 1698431365
transform 1 0 53088 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698431365
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698431365
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_37
timestamp 1698431365
transform 1 0 5488 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_47
timestamp 1698431365
transform 1 0 6608 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_51
timestamp 1698431365
transform 1 0 7056 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_54
timestamp 1698431365
transform 1 0 7392 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_74
timestamp 1698431365
transform 1 0 9632 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_78
timestamp 1698431365
transform 1 0 10080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_80
timestamp 1698431365
transform 1 0 10304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_92
timestamp 1698431365
transform 1 0 11648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_96
timestamp 1698431365
transform 1 0 12096 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_104
timestamp 1698431365
transform 1 0 12992 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698431365
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_123
timestamp 1698431365
transform 1 0 15120 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_127
timestamp 1698431365
transform 1 0 15568 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_129
timestamp 1698431365
transform 1 0 15792 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698431365
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_171
timestamp 1698431365
transform 1 0 20496 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_177
timestamp 1698431365
transform 1 0 21168 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_193
timestamp 1698431365
transform 1 0 22960 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_197
timestamp 1698431365
transform 1 0 23408 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_199
timestamp 1698431365
transform 1 0 23632 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_226
timestamp 1698431365
transform 1 0 26656 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698431365
transform 1 0 28448 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698431365
transform 1 0 28672 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698431365
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_256
timestamp 1698431365
transform 1 0 30016 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_260
timestamp 1698431365
transform 1 0 30464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_262
timestamp 1698431365
transform 1 0 30688 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_268
timestamp 1698431365
transform 1 0 31360 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_272
timestamp 1698431365
transform 1 0 31808 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_306
timestamp 1698431365
transform 1 0 35616 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_314
timestamp 1698431365
transform 1 0 36512 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_325
timestamp 1698431365
transform 1 0 37744 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_379
timestamp 1698431365
transform 1 0 43792 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_383
timestamp 1698431365
transform 1 0 44240 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_387
timestamp 1698431365
transform 1 0 44688 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_391
timestamp 1698431365
transform 1 0 45136 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_403
timestamp 1698431365
transform 1 0 46480 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_411
timestamp 1698431365
transform 1 0 47376 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_413
timestamp 1698431365
transform 1 0 47600 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_438
timestamp 1698431365
transform 1 0 50400 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_448
timestamp 1698431365
transform 1 0 51520 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_452
timestamp 1698431365
transform 1 0 51968 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_454
timestamp 1698431365
transform 1 0 52192 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_457
timestamp 1698431365
transform 1 0 52528 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_2
timestamp 1698431365
transform 1 0 1568 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_42
timestamp 1698431365
transform 1 0 6048 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_46
timestamp 1698431365
transform 1 0 6496 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_54
timestamp 1698431365
transform 1 0 7392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698431365
transform 1 0 8960 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_72
timestamp 1698431365
transform 1 0 9408 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_136
timestamp 1698431365
transform 1 0 16576 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698431365
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_150
timestamp 1698431365
transform 1 0 18144 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698431365
transform 1 0 18592 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_187
timestamp 1698431365
transform 1 0 22288 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_203
timestamp 1698431365
transform 1 0 24080 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_207
timestamp 1698431365
transform 1 0 24528 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698431365
transform 1 0 24752 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_212
timestamp 1698431365
transform 1 0 25088 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_247
timestamp 1698431365
transform 1 0 29008 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_256
timestamp 1698431365
transform 1 0 30016 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_260
timestamp 1698431365
transform 1 0 30464 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_266
timestamp 1698431365
transform 1 0 31136 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_270
timestamp 1698431365
transform 1 0 31584 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_278
timestamp 1698431365
transform 1 0 32480 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_282
timestamp 1698431365
transform 1 0 32928 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_290
timestamp 1698431365
transform 1 0 33824 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_296
timestamp 1698431365
transform 1 0 34496 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_300
timestamp 1698431365
transform 1 0 34944 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_304
timestamp 1698431365
transform 1 0 35392 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_315
timestamp 1698431365
transform 1 0 36624 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_331
timestamp 1698431365
transform 1 0 38416 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_338
timestamp 1698431365
transform 1 0 39200 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_346
timestamp 1698431365
transform 1 0 40096 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_358
timestamp 1698431365
transform 1 0 41440 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_362
timestamp 1698431365
transform 1 0 41888 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_418
timestamp 1698431365
transform 1 0 48160 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_422
timestamp 1698431365
transform 1 0 48608 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_426
timestamp 1698431365
transform 1 0 49056 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_31
timestamp 1698431365
transform 1 0 4816 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_53
timestamp 1698431365
transform 1 0 7280 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_69
timestamp 1698431365
transform 1 0 9072 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_73
timestamp 1698431365
transform 1 0 9520 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_89
timestamp 1698431365
transform 1 0 11312 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_95
timestamp 1698431365
transform 1 0 11984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_99
timestamp 1698431365
transform 1 0 12432 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_103
timestamp 1698431365
transform 1 0 12880 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_107
timestamp 1698431365
transform 1 0 13328 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_139
timestamp 1698431365
transform 1 0 16912 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_142
timestamp 1698431365
transform 1 0 17248 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_150
timestamp 1698431365
transform 1 0 18144 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_154
timestamp 1698431365
transform 1 0 18592 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_171
timestamp 1698431365
transform 1 0 20496 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_177
timestamp 1698431365
transform 1 0 21168 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_216
timestamp 1698431365
transform 1 0 25536 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_220
timestamp 1698431365
transform 1 0 25984 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_236
timestamp 1698431365
transform 1 0 27776 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_240
timestamp 1698431365
transform 1 0 28224 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_242
timestamp 1698431365
transform 1 0 28448 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_295
timestamp 1698431365
transform 1 0 34384 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_312
timestamp 1698431365
transform 1 0 36288 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_314
timestamp 1698431365
transform 1 0 36512 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698431365
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_333
timestamp 1698431365
transform 1 0 38640 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_345
timestamp 1698431365
transform 1 0 39984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_349
timestamp 1698431365
transform 1 0 40432 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_357
timestamp 1698431365
transform 1 0 41328 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_372
timestamp 1698431365
transform 1 0 43008 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_376
timestamp 1698431365
transform 1 0 43456 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_387
timestamp 1698431365
transform 1 0 44688 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_451
timestamp 1698431365
transform 1 0 51856 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_457
timestamp 1698431365
transform 1 0 52528 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_2
timestamp 1698431365
transform 1 0 1568 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_34
timestamp 1698431365
transform 1 0 5152 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_41
timestamp 1698431365
transform 1 0 5936 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_49
timestamp 1698431365
transform 1 0 6832 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_51
timestamp 1698431365
transform 1 0 7056 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_56
timestamp 1698431365
transform 1 0 7616 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_64
timestamp 1698431365
transform 1 0 8512 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_122
timestamp 1698431365
transform 1 0 15008 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_126
timestamp 1698431365
transform 1 0 15456 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_179
timestamp 1698431365
transform 1 0 21392 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698431365
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698431365
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_212
timestamp 1698431365
transform 1 0 25088 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_216
timestamp 1698431365
transform 1 0 25536 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_220
timestamp 1698431365
transform 1 0 25984 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_224
timestamp 1698431365
transform 1 0 26432 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_282
timestamp 1698431365
transform 1 0 32928 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_290
timestamp 1698431365
transform 1 0 33824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_318
timestamp 1698431365
transform 1 0 36960 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_322
timestamp 1698431365
transform 1 0 37408 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_326
timestamp 1698431365
transform 1 0 37856 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_330
timestamp 1698431365
transform 1 0 38304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_332
timestamp 1698431365
transform 1 0 38528 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_349
timestamp 1698431365
transform 1 0 40432 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_352
timestamp 1698431365
transform 1 0 40768 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_356
timestamp 1698431365
transform 1 0 41216 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_359
timestamp 1698431365
transform 1 0 41552 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_367
timestamp 1698431365
transform 1 0 42448 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_371
timestamp 1698431365
transform 1 0 42896 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_373
timestamp 1698431365
transform 1 0 43120 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_382
timestamp 1698431365
transform 1 0 44128 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_384
timestamp 1698431365
transform 1 0 44352 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_387
timestamp 1698431365
transform 1 0 44688 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_391
timestamp 1698431365
transform 1 0 45136 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_395
timestamp 1698431365
transform 1 0 45584 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_411
timestamp 1698431365
transform 1 0 47376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_415
timestamp 1698431365
transform 1 0 47824 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_417
timestamp 1698431365
transform 1 0 48048 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_428
timestamp 1698431365
transform 1 0 49280 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_444
timestamp 1698431365
transform 1 0 51072 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_452
timestamp 1698431365
transform 1 0 51968 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_456
timestamp 1698431365
transform 1 0 52416 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_2
timestamp 1698431365
transform 1 0 1568 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_6
timestamp 1698431365
transform 1 0 2016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_8
timestamp 1698431365
transform 1 0 2240 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_15
timestamp 1698431365
transform 1 0 3024 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_19
timestamp 1698431365
transform 1 0 3472 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_27
timestamp 1698431365
transform 1 0 4368 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698431365
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_45
timestamp 1698431365
transform 1 0 6384 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_53
timestamp 1698431365
transform 1 0 7280 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_63
timestamp 1698431365
transform 1 0 8400 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_71
timestamp 1698431365
transform 1 0 9296 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_81
timestamp 1698431365
transform 1 0 10416 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_85
timestamp 1698431365
transform 1 0 10864 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_92
timestamp 1698431365
transform 1 0 11648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_96
timestamp 1698431365
transform 1 0 12096 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_104
timestamp 1698431365
transform 1 0 12992 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_107
timestamp 1698431365
transform 1 0 13328 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_123
timestamp 1698431365
transform 1 0 15120 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_131
timestamp 1698431365
transform 1 0 16016 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_145
timestamp 1698431365
transform 1 0 17584 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_149
timestamp 1698431365
transform 1 0 18032 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_157
timestamp 1698431365
transform 1 0 18928 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_166
timestamp 1698431365
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_173
timestamp 1698431365
transform 1 0 20720 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_177
timestamp 1698431365
transform 1 0 21168 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_181
timestamp 1698431365
transform 1 0 21616 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_197
timestamp 1698431365
transform 1 0 23408 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_201
timestamp 1698431365
transform 1 0 23856 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_203
timestamp 1698431365
transform 1 0 24080 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_226
timestamp 1698431365
transform 1 0 26656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_230
timestamp 1698431365
transform 1 0 27104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_234
timestamp 1698431365
transform 1 0 27552 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_242
timestamp 1698431365
transform 1 0 28448 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_244
timestamp 1698431365
transform 1 0 28672 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_247
timestamp 1698431365
transform 1 0 29008 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_249
timestamp 1698431365
transform 1 0 29232 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_262
timestamp 1698431365
transform 1 0 30688 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_266
timestamp 1698431365
transform 1 0 31136 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_273
timestamp 1698431365
transform 1 0 31920 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_313
timestamp 1698431365
transform 1 0 36400 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_317
timestamp 1698431365
transform 1 0 36848 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_321
timestamp 1698431365
transform 1 0 37296 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_330
timestamp 1698431365
transform 1 0 38304 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_346
timestamp 1698431365
transform 1 0 40096 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_352
timestamp 1698431365
transform 1 0 40768 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_356
timestamp 1698431365
transform 1 0 41216 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_358
timestamp 1698431365
transform 1 0 41440 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_383
timestamp 1698431365
transform 1 0 44240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_393
timestamp 1698431365
transform 1 0 45360 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_401
timestamp 1698431365
transform 1 0 46256 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_444
timestamp 1698431365
transform 1 0 51072 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_452
timestamp 1698431365
transform 1 0 51968 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_454
timestamp 1698431365
transform 1 0 52192 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_32_457
timestamp 1698431365
transform 1 0 52528 0 1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_46
timestamp 1698431365
transform 1 0 6496 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_69
timestamp 1698431365
transform 1 0 9072 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_72
timestamp 1698431365
transform 1 0 9408 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_100
timestamp 1698431365
transform 1 0 12544 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_106
timestamp 1698431365
transform 1 0 13216 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_110
timestamp 1698431365
transform 1 0 13664 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_114
timestamp 1698431365
transform 1 0 14112 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_128
timestamp 1698431365
transform 1 0 15680 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_132
timestamp 1698431365
transform 1 0 16128 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_154
timestamp 1698431365
transform 1 0 18592 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_158
timestamp 1698431365
transform 1 0 19040 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_197
timestamp 1698431365
transform 1 0 23408 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_205
timestamp 1698431365
transform 1 0 24304 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698431365
transform 1 0 24752 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_212
timestamp 1698431365
transform 1 0 25088 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_216
timestamp 1698431365
transform 1 0 25536 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_218
timestamp 1698431365
transform 1 0 25760 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_250
timestamp 1698431365
transform 1 0 29344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_254
timestamp 1698431365
transform 1 0 29792 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_270
timestamp 1698431365
transform 1 0 31584 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_278
timestamp 1698431365
transform 1 0 32480 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_282
timestamp 1698431365
transform 1 0 32928 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_296
timestamp 1698431365
transform 1 0 34496 0 -1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_312
timestamp 1698431365
transform 1 0 36288 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_320
timestamp 1698431365
transform 1 0 37184 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_324
timestamp 1698431365
transform 1 0 37632 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_344
timestamp 1698431365
transform 1 0 39872 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_352
timestamp 1698431365
transform 1 0 40768 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_354
timestamp 1698431365
transform 1 0 40992 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_371
timestamp 1698431365
transform 1 0 42896 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_379
timestamp 1698431365
transform 1 0 43792 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_410
timestamp 1698431365
transform 1 0 47264 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_418
timestamp 1698431365
transform 1 0 48160 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_33_422
timestamp 1698431365
transform 1 0 48608 0 -1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_430
timestamp 1698431365
transform 1 0 49504 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_434
timestamp 1698431365
transform 1 0 49952 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_2
timestamp 1698431365
transform 1 0 1568 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_18
timestamp 1698431365
transform 1 0 3360 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_26
timestamp 1698431365
transform 1 0 4256 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_30
timestamp 1698431365
transform 1 0 4704 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_33
timestamp 1698431365
transform 1 0 5040 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_37
timestamp 1698431365
transform 1 0 5488 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_69
timestamp 1698431365
transform 1 0 9072 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_104
timestamp 1698431365
transform 1 0 12992 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_113
timestamp 1698431365
transform 1 0 14000 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_129
timestamp 1698431365
transform 1 0 15792 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_141
timestamp 1698431365
transform 1 0 17136 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_157
timestamp 1698431365
transform 1 0 18928 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_165
timestamp 1698431365
transform 1 0 19824 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_169
timestamp 1698431365
transform 1 0 20272 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_185
timestamp 1698431365
transform 1 0 22064 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_193
timestamp 1698431365
transform 1 0 22960 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_204
timestamp 1698431365
transform 1 0 24192 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_208
timestamp 1698431365
transform 1 0 24640 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_210
timestamp 1698431365
transform 1 0 24864 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_219
timestamp 1698431365
transform 1 0 25872 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_223
timestamp 1698431365
transform 1 0 26320 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_239
timestamp 1698431365
transform 1 0 28112 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_243
timestamp 1698431365
transform 1 0 28560 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_247
timestamp 1698431365
transform 1 0 29008 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_249
timestamp 1698431365
transform 1 0 29232 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_269
timestamp 1698431365
transform 1 0 31472 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_273
timestamp 1698431365
transform 1 0 31920 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_281
timestamp 1698431365
transform 1 0 32816 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_285
timestamp 1698431365
transform 1 0 33264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_310
timestamp 1698431365
transform 1 0 36064 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_314
timestamp 1698431365
transform 1 0 36512 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_325
timestamp 1698431365
transform 1 0 37744 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_331
timestamp 1698431365
transform 1 0 38416 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_347
timestamp 1698431365
transform 1 0 40208 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_351
timestamp 1698431365
transform 1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_353
timestamp 1698431365
transform 1 0 40880 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_360
timestamp 1698431365
transform 1 0 41664 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_370
timestamp 1698431365
transform 1 0 42784 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_378
timestamp 1698431365
transform 1 0 43680 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_382
timestamp 1698431365
transform 1 0 44128 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_384
timestamp 1698431365
transform 1 0 44352 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_387
timestamp 1698431365
transform 1 0 44688 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_34_419
timestamp 1698431365
transform 1 0 48272 0 1 29792
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_34_441
timestamp 1698431365
transform 1 0 50736 0 1 29792
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_449
timestamp 1698431365
transform 1 0 51632 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_34_457
timestamp 1698431365
transform 1 0 52528 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_2
timestamp 1698431365
transform 1 0 1568 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_34
timestamp 1698431365
transform 1 0 5152 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_42
timestamp 1698431365
transform 1 0 6048 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_57
timestamp 1698431365
transform 1 0 7728 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_65
timestamp 1698431365
transform 1 0 8624 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_69
timestamp 1698431365
transform 1 0 9072 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_84
timestamp 1698431365
transform 1 0 10752 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_86
timestamp 1698431365
transform 1 0 10976 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_116
timestamp 1698431365
transform 1 0 14336 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_120
timestamp 1698431365
transform 1 0 14784 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_122
timestamp 1698431365
transform 1 0 15008 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_135
timestamp 1698431365
transform 1 0 16464 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_139
timestamp 1698431365
transform 1 0 16912 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_142
timestamp 1698431365
transform 1 0 17248 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_35_156
timestamp 1698431365
transform 1 0 18816 0 -1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_188
timestamp 1698431365
transform 1 0 22400 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_204
timestamp 1698431365
transform 1 0 24192 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_222
timestamp 1698431365
transform 1 0 26208 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_226
timestamp 1698431365
transform 1 0 26656 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_242
timestamp 1698431365
transform 1 0 28448 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_246
timestamp 1698431365
transform 1 0 28896 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_248
timestamp 1698431365
transform 1 0 29120 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_282
timestamp 1698431365
transform 1 0 32928 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_286
timestamp 1698431365
transform 1 0 33376 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_304
timestamp 1698431365
transform 1 0 35392 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_308
timestamp 1698431365
transform 1 0 35840 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_319
timestamp 1698431365
transform 1 0 37072 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_321
timestamp 1698431365
transform 1 0 37296 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_35_341
timestamp 1698431365
transform 1 0 39536 0 -1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_349
timestamp 1698431365
transform 1 0 40432 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_352
timestamp 1698431365
transform 1 0 40768 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_368
timestamp 1698431365
transform 1 0 42560 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_35_391
timestamp 1698431365
transform 1 0 45136 0 -1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_407
timestamp 1698431365
transform 1 0 46928 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_411
timestamp 1698431365
transform 1 0 47376 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_413
timestamp 1698431365
transform 1 0 47600 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_432
timestamp 1698431365
transform 1 0 49728 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_2
timestamp 1698431365
transform 1 0 1568 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_18
timestamp 1698431365
transform 1 0 3360 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_26
timestamp 1698431365
transform 1 0 4256 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_30
timestamp 1698431365
transform 1 0 4704 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_33
timestamp 1698431365
transform 1 0 5040 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_53
timestamp 1698431365
transform 1 0 7280 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_61
timestamp 1698431365
transform 1 0 8176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_79
timestamp 1698431365
transform 1 0 10192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_85
timestamp 1698431365
transform 1 0 10864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_89
timestamp 1698431365
transform 1 0 11312 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_107
timestamp 1698431365
transform 1 0 13328 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_115
timestamp 1698431365
transform 1 0 14224 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_117
timestamp 1698431365
transform 1 0 14448 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_120
timestamp 1698431365
transform 1 0 14784 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_136
timestamp 1698431365
transform 1 0 16576 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_140
timestamp 1698431365
transform 1 0 17024 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_167
timestamp 1698431365
transform 1 0 20048 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698431365
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_177
timestamp 1698431365
transform 1 0 21168 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_193
timestamp 1698431365
transform 1 0 22960 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_210
timestamp 1698431365
transform 1 0 24864 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_247
timestamp 1698431365
transform 1 0 29008 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_36_251
timestamp 1698431365
transform 1 0 29456 0 1 31360
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_267
timestamp 1698431365
transform 1 0 31248 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_271
timestamp 1698431365
transform 1 0 31696 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_275
timestamp 1698431365
transform 1 0 32144 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_283
timestamp 1698431365
transform 1 0 33040 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_287
timestamp 1698431365
transform 1 0 33488 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_291
timestamp 1698431365
transform 1 0 33936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_300
timestamp 1698431365
transform 1 0 34944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_304
timestamp 1698431365
transform 1 0 35392 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_312
timestamp 1698431365
transform 1 0 36288 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_314
timestamp 1698431365
transform 1 0 36512 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_317
timestamp 1698431365
transform 1 0 36848 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_321
timestamp 1698431365
transform 1 0 37296 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_325
timestamp 1698431365
transform 1 0 37744 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_333
timestamp 1698431365
transform 1 0 38640 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_339
timestamp 1698431365
transform 1 0 39312 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_349
timestamp 1698431365
transform 1 0 40432 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_358
timestamp 1698431365
transform 1 0 41440 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_362
timestamp 1698431365
transform 1 0 41888 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_364
timestamp 1698431365
transform 1 0 42112 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_383
timestamp 1698431365
transform 1 0 44240 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_416
timestamp 1698431365
transform 1 0 47936 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_420
timestamp 1698431365
transform 1 0 48384 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_428
timestamp 1698431365
transform 1 0 49280 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_432
timestamp 1698431365
transform 1 0 49728 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_448
timestamp 1698431365
transform 1 0 51520 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_36_452
timestamp 1698431365
transform 1 0 51968 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_454
timestamp 1698431365
transform 1 0 52192 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_36_457
timestamp 1698431365
transform 1 0 52528 0 1 31360
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_31
timestamp 1698431365
transform 1 0 4816 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_33
timestamp 1698431365
transform 1 0 5040 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_49
timestamp 1698431365
transform 1 0 6832 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_53
timestamp 1698431365
transform 1 0 7280 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_69
timestamp 1698431365
transform 1 0 9072 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_77
timestamp 1698431365
transform 1 0 9968 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_93
timestamp 1698431365
transform 1 0 11760 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_101
timestamp 1698431365
transform 1 0 12656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_103
timestamp 1698431365
transform 1 0 12880 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_118
timestamp 1698431365
transform 1 0 14560 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_129
timestamp 1698431365
transform 1 0 15792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_135
timestamp 1698431365
transform 1 0 16464 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_137
timestamp 1698431365
transform 1 0 16688 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_142
timestamp 1698431365
transform 1 0 17248 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_179
timestamp 1698431365
transform 1 0 21392 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_183
timestamp 1698431365
transform 1 0 21840 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_196
timestamp 1698431365
transform 1 0 23296 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_200
timestamp 1698431365
transform 1 0 23744 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_212
timestamp 1698431365
transform 1 0 25088 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_220
timestamp 1698431365
transform 1 0 25984 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_224
timestamp 1698431365
transform 1 0 26432 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_240
timestamp 1698431365
transform 1 0 28224 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_248
timestamp 1698431365
transform 1 0 29120 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_252
timestamp 1698431365
transform 1 0 29568 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_254
timestamp 1698431365
transform 1 0 29792 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_267
timestamp 1698431365
transform 1 0 31248 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_271
timestamp 1698431365
transform 1 0 31696 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_282
timestamp 1698431365
transform 1 0 32928 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_284
timestamp 1698431365
transform 1 0 33152 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_332
timestamp 1698431365
transform 1 0 38528 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_336
timestamp 1698431365
transform 1 0 38976 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698431365
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_358
timestamp 1698431365
transform 1 0 41440 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_366
timestamp 1698431365
transform 1 0 42336 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_37_379
timestamp 1698431365
transform 1 0 43792 0 -1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_37_411
timestamp 1698431365
transform 1 0 47376 0 -1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_419
timestamp 1698431365
transform 1 0 48272 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_37_422
timestamp 1698431365
transform 1 0 48608 0 -1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_438
timestamp 1698431365
transform 1 0 50400 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698431365
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698431365
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_48
timestamp 1698431365
transform 1 0 6720 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_56
timestamp 1698431365
transform 1 0 7616 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_64
timestamp 1698431365
transform 1 0 8512 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_68
timestamp 1698431365
transform 1 0 8960 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_75
timestamp 1698431365
transform 1 0 9744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_90
timestamp 1698431365
transform 1 0 11424 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_94
timestamp 1698431365
transform 1 0 11872 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_102
timestamp 1698431365
transform 1 0 12768 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_104
timestamp 1698431365
transform 1 0 12992 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_107
timestamp 1698431365
transform 1 0 13328 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_111
timestamp 1698431365
transform 1 0 13776 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_113
timestamp 1698431365
transform 1 0 14000 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_164
timestamp 1698431365
transform 1 0 19712 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_168
timestamp 1698431365
transform 1 0 20160 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_185
timestamp 1698431365
transform 1 0 22064 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_193
timestamp 1698431365
transform 1 0 22960 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_200
timestamp 1698431365
transform 1 0 23744 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_204
timestamp 1698431365
transform 1 0 24192 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_212
timestamp 1698431365
transform 1 0 25088 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_214
timestamp 1698431365
transform 1 0 25312 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_220
timestamp 1698431365
transform 1 0 25984 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_224
timestamp 1698431365
transform 1 0 26432 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_240
timestamp 1698431365
transform 1 0 28224 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_244
timestamp 1698431365
transform 1 0 28672 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_247
timestamp 1698431365
transform 1 0 29008 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_249
timestamp 1698431365
transform 1 0 29232 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_269
timestamp 1698431365
transform 1 0 31472 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_277
timestamp 1698431365
transform 1 0 32368 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_279
timestamp 1698431365
transform 1 0 32592 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_292
timestamp 1698431365
transform 1 0 34048 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_296
timestamp 1698431365
transform 1 0 34496 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_312
timestamp 1698431365
transform 1 0 36288 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_314
timestamp 1698431365
transform 1 0 36512 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698431365
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_349
timestamp 1698431365
transform 1 0 40432 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_352
timestamp 1698431365
transform 1 0 40768 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_362
timestamp 1698431365
transform 1 0 41888 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_378
timestamp 1698431365
transform 1 0 43680 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_382
timestamp 1698431365
transform 1 0 44128 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_384
timestamp 1698431365
transform 1 0 44352 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_387
timestamp 1698431365
transform 1 0 44688 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_391
timestamp 1698431365
transform 1 0 45136 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_38_400
timestamp 1698431365
transform 1 0 46144 0 1 32928
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_416
timestamp 1698431365
transform 1 0 47936 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_422
timestamp 1698431365
transform 1 0 48608 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_430
timestamp 1698431365
transform 1 0 49504 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_432
timestamp 1698431365
transform 1 0 49728 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_441
timestamp 1698431365
transform 1 0 50736 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_449
timestamp 1698431365
transform 1 0 51632 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_38_453
timestamp 1698431365
transform 1 0 52080 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_38_457
timestamp 1698431365
transform 1 0 52528 0 1 32928
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_2
timestamp 1698431365
transform 1 0 1568 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_18
timestamp 1698431365
transform 1 0 3360 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_26
timestamp 1698431365
transform 1 0 4256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_30
timestamp 1698431365
transform 1 0 4704 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_38
timestamp 1698431365
transform 1 0 5600 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_47
timestamp 1698431365
transform 1 0 6608 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_63
timestamp 1698431365
transform 1 0 8400 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_67
timestamp 1698431365
transform 1 0 8848 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_69
timestamp 1698431365
transform 1 0 9072 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_72
timestamp 1698431365
transform 1 0 9408 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_109
timestamp 1698431365
transform 1 0 13552 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_113
timestamp 1698431365
transform 1 0 14000 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_121
timestamp 1698431365
transform 1 0 14896 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_125
timestamp 1698431365
transform 1 0 15344 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_128
timestamp 1698431365
transform 1 0 15680 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698431365
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_142
timestamp 1698431365
transform 1 0 17248 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_152
timestamp 1698431365
transform 1 0 18368 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_154
timestamp 1698431365
transform 1 0 18592 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_157
timestamp 1698431365
transform 1 0 18928 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_161
timestamp 1698431365
transform 1 0 19376 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_198
timestamp 1698431365
transform 1 0 23520 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_206
timestamp 1698431365
transform 1 0 24416 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_212
timestamp 1698431365
transform 1 0 25088 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_214
timestamp 1698431365
transform 1 0 25312 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_39_223
timestamp 1698431365
transform 1 0 26320 0 -1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_239
timestamp 1698431365
transform 1 0 28112 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_243
timestamp 1698431365
transform 1 0 28560 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_246
timestamp 1698431365
transform 1 0 28896 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_254
timestamp 1698431365
transform 1 0 29792 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_256
timestamp 1698431365
transform 1 0 30016 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_262
timestamp 1698431365
transform 1 0 30688 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_266
timestamp 1698431365
transform 1 0 31136 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_274
timestamp 1698431365
transform 1 0 32032 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_278
timestamp 1698431365
transform 1 0 32480 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_39_282
timestamp 1698431365
transform 1 0 32928 0 -1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_314
timestamp 1698431365
transform 1 0 36512 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_317
timestamp 1698431365
transform 1 0 36848 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_325
timestamp 1698431365
transform 1 0 37744 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_327
timestamp 1698431365
transform 1 0 37968 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_339
timestamp 1698431365
transform 1 0 39312 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_346
timestamp 1698431365
transform 1 0 40096 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_360
timestamp 1698431365
transform 1 0 41664 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_362
timestamp 1698431365
transform 1 0 41888 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_39_382
timestamp 1698431365
transform 1 0 44128 0 -1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_390
timestamp 1698431365
transform 1 0 45024 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_45
timestamp 1698431365
transform 1 0 6384 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_53
timestamp 1698431365
transform 1 0 7280 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_57
timestamp 1698431365
transform 1 0 7728 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_59
timestamp 1698431365
transform 1 0 7952 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_62
timestamp 1698431365
transform 1 0 8288 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_77
timestamp 1698431365
transform 1 0 9968 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_93
timestamp 1698431365
transform 1 0 11760 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698431365
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_107
timestamp 1698431365
transform 1 0 13328 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_111
timestamp 1698431365
transform 1 0 13776 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_124
timestamp 1698431365
transform 1 0 15232 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_128
timestamp 1698431365
transform 1 0 15680 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_144
timestamp 1698431365
transform 1 0 17472 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_146
timestamp 1698431365
transform 1 0 17696 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_159
timestamp 1698431365
transform 1 0 19152 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_163
timestamp 1698431365
transform 1 0 19600 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698431365
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_177
timestamp 1698431365
transform 1 0 21168 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_193
timestamp 1698431365
transform 1 0 22960 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_201
timestamp 1698431365
transform 1 0 23856 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_203
timestamp 1698431365
transform 1 0 24080 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_211
timestamp 1698431365
transform 1 0 24976 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_244
timestamp 1698431365
transform 1 0 28672 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_278
timestamp 1698431365
transform 1 0 32480 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_282
timestamp 1698431365
transform 1 0 32928 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_298
timestamp 1698431365
transform 1 0 34720 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_306
timestamp 1698431365
transform 1 0 35616 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_309
timestamp 1698431365
transform 1 0 35952 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_313
timestamp 1698431365
transform 1 0 36400 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_342
timestamp 1698431365
transform 1 0 39648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_364
timestamp 1698431365
transform 1 0 42112 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_371
timestamp 1698431365
transform 1 0 42896 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_375
timestamp 1698431365
transform 1 0 43344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_382
timestamp 1698431365
transform 1 0 44128 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_384
timestamp 1698431365
transform 1 0 44352 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_392
timestamp 1698431365
transform 1 0 45248 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_424
timestamp 1698431365
transform 1 0 48832 0 1 34496
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_440
timestamp 1698431365
transform 1 0 50624 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_448
timestamp 1698431365
transform 1 0 51520 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_40_452
timestamp 1698431365
transform 1 0 51968 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_454
timestamp 1698431365
transform 1 0 52192 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_457
timestamp 1698431365
transform 1 0 52528 0 1 34496
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_2
timestamp 1698431365
transform 1 0 1568 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_18
timestamp 1698431365
transform 1 0 3360 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_26
timestamp 1698431365
transform 1 0 4256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_30
timestamp 1698431365
transform 1 0 4704 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_33
timestamp 1698431365
transform 1 0 5040 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_40
timestamp 1698431365
transform 1 0 5824 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_48
timestamp 1698431365
transform 1 0 6720 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_52
timestamp 1698431365
transform 1 0 7168 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_72
timestamp 1698431365
transform 1 0 9408 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_41_104
timestamp 1698431365
transform 1 0 12992 0 -1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_120
timestamp 1698431365
transform 1 0 14784 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_41_142
timestamp 1698431365
transform 1 0 17248 0 -1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_174
timestamp 1698431365
transform 1 0 20832 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_182
timestamp 1698431365
transform 1 0 21728 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_198
timestamp 1698431365
transform 1 0 23520 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_202
timestamp 1698431365
transform 1 0 23968 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698431365
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698431365
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_338
timestamp 1698431365
transform 1 0 39200 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_346
timestamp 1698431365
transform 1 0 40096 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_352
timestamp 1698431365
transform 1 0 40768 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_356
timestamp 1698431365
transform 1 0 41216 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_360
timestamp 1698431365
transform 1 0 41664 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_364
timestamp 1698431365
transform 1 0 42112 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_394
timestamp 1698431365
transform 1 0 45472 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_41_406
timestamp 1698431365
transform 1 0 46816 0 -1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_414
timestamp 1698431365
transform 1 0 47712 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_418
timestamp 1698431365
transform 1 0 48160 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_422
timestamp 1698431365
transform 1 0 48608 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_434
timestamp 1698431365
transform 1 0 49952 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_438
timestamp 1698431365
transform 1 0 50400 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_2
timestamp 1698431365
transform 1 0 1568 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_18
timestamp 1698431365
transform 1 0 3360 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_26
timestamp 1698431365
transform 1 0 4256 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_30
timestamp 1698431365
transform 1 0 4704 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_33
timestamp 1698431365
transform 1 0 5040 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_37
timestamp 1698431365
transform 1 0 5488 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_44
timestamp 1698431365
transform 1 0 6272 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_60
timestamp 1698431365
transform 1 0 8064 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_74
timestamp 1698431365
transform 1 0 9632 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_82
timestamp 1698431365
transform 1 0 10528 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_84
timestamp 1698431365
transform 1 0 10752 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_87
timestamp 1698431365
transform 1 0 11088 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_103
timestamp 1698431365
transform 1 0 12880 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_107
timestamp 1698431365
transform 1 0 13328 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_115
timestamp 1698431365
transform 1 0 14224 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_129
timestamp 1698431365
transform 1 0 15792 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_133
timestamp 1698431365
transform 1 0 16240 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_141
timestamp 1698431365
transform 1 0 17136 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_166
timestamp 1698431365
transform 1 0 19936 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_170
timestamp 1698431365
transform 1 0 20384 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_174
timestamp 1698431365
transform 1 0 20832 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_177
timestamp 1698431365
transform 1 0 21168 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_179
timestamp 1698431365
transform 1 0 21392 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_211
timestamp 1698431365
transform 1 0 24976 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_227
timestamp 1698431365
transform 1 0 26768 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_231
timestamp 1698431365
transform 1 0 27216 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_247
timestamp 1698431365
transform 1 0 29008 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_251
timestamp 1698431365
transform 1 0 29456 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_255
timestamp 1698431365
transform 1 0 29904 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_287
timestamp 1698431365
transform 1 0 33488 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_291
timestamp 1698431365
transform 1 0 33936 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_309
timestamp 1698431365
transform 1 0 35952 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_313
timestamp 1698431365
transform 1 0 36400 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_317
timestamp 1698431365
transform 1 0 36848 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_321
timestamp 1698431365
transform 1 0 37296 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_329
timestamp 1698431365
transform 1 0 38192 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_341
timestamp 1698431365
transform 1 0 39536 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_345
timestamp 1698431365
transform 1 0 39984 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_377
timestamp 1698431365
transform 1 0 43568 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_387
timestamp 1698431365
transform 1 0 44688 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_395
timestamp 1698431365
transform 1 0 45584 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_397
timestamp 1698431365
transform 1 0 45808 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_427
timestamp 1698431365
transform 1 0 49168 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_449
timestamp 1698431365
transform 1 0 51632 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_453
timestamp 1698431365
transform 1 0 52080 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_457
timestamp 1698431365
transform 1 0 52528 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_47
timestamp 1698431365
transform 1 0 6608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_57
timestamp 1698431365
transform 1 0 7728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_61
timestamp 1698431365
transform 1 0 8176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_114
timestamp 1698431365
transform 1 0 14112 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_118
timestamp 1698431365
transform 1 0 14560 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_132
timestamp 1698431365
transform 1 0 16128 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698431365
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698431365
transform 1 0 17248 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_150
timestamp 1698431365
transform 1 0 18144 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_164
timestamp 1698431365
transform 1 0 19712 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_168
timestamp 1698431365
transform 1 0 20160 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_200
timestamp 1698431365
transform 1 0 23744 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_208
timestamp 1698431365
transform 1 0 24640 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_224
timestamp 1698431365
transform 1 0 26432 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_228
timestamp 1698431365
transform 1 0 26880 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_254
timestamp 1698431365
transform 1 0 29792 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698431365
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698431365
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_282
timestamp 1698431365
transform 1 0 32928 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_298
timestamp 1698431365
transform 1 0 34720 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_306
timestamp 1698431365
transform 1 0 35616 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_310
timestamp 1698431365
transform 1 0 36064 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_312
timestamp 1698431365
transform 1 0 36288 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_315
timestamp 1698431365
transform 1 0 36624 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_352
timestamp 1698431365
transform 1 0 40768 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_368
timestamp 1698431365
transform 1 0 42560 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_384
timestamp 1698431365
transform 1 0 44352 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_416
timestamp 1698431365
transform 1 0 47936 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_430
timestamp 1698431365
transform 1 0 49504 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_434
timestamp 1698431365
transform 1 0 49952 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_2
timestamp 1698431365
transform 1 0 1568 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_18
timestamp 1698431365
transform 1 0 3360 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_26
timestamp 1698431365
transform 1 0 4256 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_37
timestamp 1698431365
transform 1 0 5488 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_44
timestamp 1698431365
transform 1 0 6272 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_60
timestamp 1698431365
transform 1 0 8064 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_68
timestamp 1698431365
transform 1 0 8960 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_77
timestamp 1698431365
transform 1 0 9968 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_93
timestamp 1698431365
transform 1 0 11760 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_101
timestamp 1698431365
transform 1 0 12656 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_107
timestamp 1698431365
transform 1 0 13328 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_139
timestamp 1698431365
transform 1 0 16912 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_177
timestamp 1698431365
transform 1 0 21168 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_181
timestamp 1698431365
transform 1 0 21616 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_213
timestamp 1698431365
transform 1 0 25200 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_226
timestamp 1698431365
transform 1 0 26656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_230
timestamp 1698431365
transform 1 0 27104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_232
timestamp 1698431365
transform 1 0 27328 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_247
timestamp 1698431365
transform 1 0 29008 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_251
timestamp 1698431365
transform 1 0 29456 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_255
timestamp 1698431365
transform 1 0 29904 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_270
timestamp 1698431365
transform 1 0 31584 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_277
timestamp 1698431365
transform 1 0 32368 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_281
timestamp 1698431365
transform 1 0 32816 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_284
timestamp 1698431365
transform 1 0 33152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_325
timestamp 1698431365
transform 1 0 37744 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_329
timestamp 1698431365
transform 1 0 38192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_331
timestamp 1698431365
transform 1 0 38416 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_337
timestamp 1698431365
transform 1 0 39088 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_345
timestamp 1698431365
transform 1 0 39984 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_349
timestamp 1698431365
transform 1 0 40432 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_351
timestamp 1698431365
transform 1 0 40656 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_358
timestamp 1698431365
transform 1 0 41440 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_374
timestamp 1698431365
transform 1 0 43232 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_382
timestamp 1698431365
transform 1 0 44128 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_413
timestamp 1698431365
transform 1 0 47600 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_445
timestamp 1698431365
transform 1 0 51184 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_453
timestamp 1698431365
transform 1 0 52080 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_457
timestamp 1698431365
transform 1 0 52528 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_2
timestamp 1698431365
transform 1 0 1568 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_34
timestamp 1698431365
transform 1 0 5152 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_50
timestamp 1698431365
transform 1 0 6944 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_67
timestamp 1698431365
transform 1 0 8848 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_69
timestamp 1698431365
transform 1 0 9072 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_72
timestamp 1698431365
transform 1 0 9408 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_79
timestamp 1698431365
transform 1 0 10192 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_95
timestamp 1698431365
transform 1 0 11984 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_103
timestamp 1698431365
transform 1 0 12880 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_106
timestamp 1698431365
transform 1 0 13216 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_122
timestamp 1698431365
transform 1 0 15008 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_126
timestamp 1698431365
transform 1 0 15456 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_142
timestamp 1698431365
transform 1 0 17248 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_146
timestamp 1698431365
transform 1 0 17696 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_150
timestamp 1698431365
transform 1 0 18144 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_158
timestamp 1698431365
transform 1 0 19040 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_45_212
timestamp 1698431365
transform 1 0 25088 0 -1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_244
timestamp 1698431365
transform 1 0 28672 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_282
timestamp 1698431365
transform 1 0 32928 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_296
timestamp 1698431365
transform 1 0 34496 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_298
timestamp 1698431365
transform 1 0 34720 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_327
timestamp 1698431365
transform 1 0 37968 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_343
timestamp 1698431365
transform 1 0 39760 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_347
timestamp 1698431365
transform 1 0 40208 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_349
timestamp 1698431365
transform 1 0 40432 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_45_352
timestamp 1698431365
transform 1 0 40768 0 -1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_45_368
timestamp 1698431365
transform 1 0 42560 0 -1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_398
timestamp 1698431365
transform 1 0 45920 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_412
timestamp 1698431365
transform 1 0 47488 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_45_422
timestamp 1698431365
transform 1 0 48608 0 -1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_45_430
timestamp 1698431365
transform 1 0 49504 0 -1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_45_434
timestamp 1698431365
transform 1 0 49952 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_2
timestamp 1698431365
transform 1 0 1568 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_18
timestamp 1698431365
transform 1 0 3360 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_26
timestamp 1698431365
transform 1 0 4256 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_30
timestamp 1698431365
transform 1 0 4704 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_49
timestamp 1698431365
transform 1 0 6832 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_57
timestamp 1698431365
transform 1 0 7728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_66
timestamp 1698431365
transform 1 0 8736 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_104
timestamp 1698431365
transform 1 0 12992 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_148
timestamp 1698431365
transform 1 0 17920 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_150
timestamp 1698431365
transform 1 0 18144 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_163
timestamp 1698431365
transform 1 0 19600 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_171
timestamp 1698431365
transform 1 0 20496 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_177
timestamp 1698431365
transform 1 0 21168 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_193
timestamp 1698431365
transform 1 0 22960 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_203
timestamp 1698431365
transform 1 0 24080 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_235
timestamp 1698431365
transform 1 0 27664 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_244
timestamp 1698431365
transform 1 0 28672 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_46_247
timestamp 1698431365
transform 1 0 29008 0 1 39200
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_279
timestamp 1698431365
transform 1 0 32592 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_295
timestamp 1698431365
transform 1 0 34384 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_46_303
timestamp 1698431365
transform 1 0 35280 0 1 39200
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_307
timestamp 1698431365
transform 1 0 35728 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_309
timestamp 1698431365
transform 1 0 35952 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_322
timestamp 1698431365
transform 1 0 37408 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_359
timestamp 1698431365
transform 1 0 41552 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_46_363
timestamp 1698431365
transform 1 0 42000 0 1 39200
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_379
timestamp 1698431365
transform 1 0 43792 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_395
timestamp 1698431365
transform 1 0 45584 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_397
timestamp 1698431365
transform 1 0 45808 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_46_403
timestamp 1698431365
transform 1 0 46480 0 1 39200
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_433
timestamp 1698431365
transform 1 0 49840 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_46_451
timestamp 1698431365
transform 1 0 51856 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_46_457
timestamp 1698431365
transform 1 0 52528 0 1 39200
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_2
timestamp 1698431365
transform 1 0 1568 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_34
timestamp 1698431365
transform 1 0 5152 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_43
timestamp 1698431365
transform 1 0 6160 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_51
timestamp 1698431365
transform 1 0 7056 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_55
timestamp 1698431365
transform 1 0 7504 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_57
timestamp 1698431365
transform 1 0 7728 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_64
timestamp 1698431365
transform 1 0 8512 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_68
timestamp 1698431365
transform 1 0 8960 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_47_72
timestamp 1698431365
transform 1 0 9408 0 -1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_104
timestamp 1698431365
transform 1 0 12992 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_120
timestamp 1698431365
transform 1 0 14784 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_128
timestamp 1698431365
transform 1 0 15680 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_138
timestamp 1698431365
transform 1 0 16800 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_142
timestamp 1698431365
transform 1 0 17248 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_150
timestamp 1698431365
transform 1 0 18144 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_185
timestamp 1698431365
transform 1 0 22064 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_189
timestamp 1698431365
transform 1 0 22512 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_208
timestamp 1698431365
transform 1 0 24640 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_212
timestamp 1698431365
transform 1 0 25088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_216
timestamp 1698431365
transform 1 0 25536 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_246
timestamp 1698431365
transform 1 0 28896 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_250
timestamp 1698431365
transform 1 0 29344 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_266
timestamp 1698431365
transform 1 0 31136 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_279
timestamp 1698431365
transform 1 0 32592 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_282
timestamp 1698431365
transform 1 0 32928 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_286
timestamp 1698431365
transform 1 0 33376 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_330
timestamp 1698431365
transform 1 0 38304 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_47_337
timestamp 1698431365
transform 1 0 39088 0 -1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_341
timestamp 1698431365
transform 1 0 39536 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_343
timestamp 1698431365
transform 1 0 39760 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_349
timestamp 1698431365
transform 1 0 40432 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_360
timestamp 1698431365
transform 1 0 41664 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_368
timestamp 1698431365
transform 1 0 42560 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_376
timestamp 1698431365
transform 1 0 43456 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_47_410
timestamp 1698431365
transform 1 0 47264 0 -1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_47_418
timestamp 1698431365
transform 1 0 48160 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_47_422
timestamp 1698431365
transform 1 0 48608 0 -1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_47_438
timestamp 1698431365
transform 1 0 50400 0 -1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_48_2
timestamp 1698431365
transform 1 0 1568 0 1 40768
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_34
timestamp 1698431365
transform 1 0 5152 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_48_37
timestamp 1698431365
transform 1 0 5488 0 1 40768
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_101
timestamp 1698431365
transform 1 0 12656 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_107
timestamp 1698431365
transform 1 0 13328 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_125
timestamp 1698431365
transform 1 0 15344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_129
timestamp 1698431365
transform 1 0 15792 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_131
timestamp 1698431365
transform 1 0 16016 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_161
timestamp 1698431365
transform 1 0 19376 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_165
timestamp 1698431365
transform 1 0 19824 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_173
timestamp 1698431365
transform 1 0 20720 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_177
timestamp 1698431365
transform 1 0 21168 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_181
timestamp 1698431365
transform 1 0 21616 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_183
timestamp 1698431365
transform 1 0 21840 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_230
timestamp 1698431365
transform 1 0 27104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_234
timestamp 1698431365
transform 1 0 27552 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_242
timestamp 1698431365
transform 1 0 28448 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_244
timestamp 1698431365
transform 1 0 28672 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_247
timestamp 1698431365
transform 1 0 29008 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_263
timestamp 1698431365
transform 1 0 30800 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_271
timestamp 1698431365
transform 1 0 31696 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_275
timestamp 1698431365
transform 1 0 32144 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_279
timestamp 1698431365
transform 1 0 32592 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_283
timestamp 1698431365
transform 1 0 33040 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_285
timestamp 1698431365
transform 1 0 33264 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_325
timestamp 1698431365
transform 1 0 37744 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_341
timestamp 1698431365
transform 1 0 39536 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_349
timestamp 1698431365
transform 1 0 40432 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_352
timestamp 1698431365
transform 1 0 40768 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_362
timestamp 1698431365
transform 1 0 41888 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_378
timestamp 1698431365
transform 1 0 43680 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_48_382
timestamp 1698431365
transform 1 0 44128 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_48_384
timestamp 1698431365
transform 1 0 44352 0 1 40768
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_387
timestamp 1698431365
transform 1 0 44688 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_48_399
timestamp 1698431365
transform 1 0 46032 0 1 40768
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_48_415
timestamp 1698431365
transform 1 0 47824 0 1 40768
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_48_457
timestamp 1698431365
transform 1 0 52528 0 1 40768
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_2
timestamp 1698431365
transform 1 0 1568 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_18
timestamp 1698431365
transform 1 0 3360 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_26
timestamp 1698431365
transform 1 0 4256 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_30
timestamp 1698431365
transform 1 0 4704 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_60
timestamp 1698431365
transform 1 0 8064 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_64
timestamp 1698431365
transform 1 0 8512 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_68
timestamp 1698431365
transform 1 0 8960 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_72
timestamp 1698431365
transform 1 0 9408 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_88
timestamp 1698431365
transform 1 0 11200 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_96
timestamp 1698431365
transform 1 0 12096 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_103
timestamp 1698431365
transform 1 0 12880 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_111
timestamp 1698431365
transform 1 0 13776 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_125
timestamp 1698431365
transform 1 0 15344 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_133
timestamp 1698431365
transform 1 0 16240 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_137
timestamp 1698431365
transform 1 0 16688 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_139
timestamp 1698431365
transform 1 0 16912 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_49_142
timestamp 1698431365
transform 1 0 17248 0 -1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_174
timestamp 1698431365
transform 1 0 20832 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_190
timestamp 1698431365
transform 1 0 22624 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_192
timestamp 1698431365
transform 1 0 22848 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_208
timestamp 1698431365
transform 1 0 24640 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_212
timestamp 1698431365
transform 1 0 25088 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_234
timestamp 1698431365
transform 1 0 27552 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_242
timestamp 1698431365
transform 1 0 28448 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_277
timestamp 1698431365
transform 1 0 32368 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_279
timestamp 1698431365
transform 1 0 32592 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_49_290
timestamp 1698431365
transform 1 0 33824 0 -1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_306
timestamp 1698431365
transform 1 0 35616 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_314
timestamp 1698431365
transform 1 0 36512 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_317
timestamp 1698431365
transform 1 0 36848 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_325
timestamp 1698431365
transform 1 0 37744 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_334
timestamp 1698431365
transform 1 0 38752 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_49_342
timestamp 1698431365
transform 1 0 39648 0 -1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_348
timestamp 1698431365
transform 1 0 40320 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_358
timestamp 1698431365
transform 1 0 41440 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_366
timestamp 1698431365
transform 1 0 42336 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_370
timestamp 1698431365
transform 1 0 42784 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_49_377
timestamp 1698431365
transform 1 0 43568 0 -1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_49_385
timestamp 1698431365
transform 1 0 44464 0 -1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_389
timestamp 1698431365
transform 1 0 44912 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_422
timestamp 1698431365
transform 1 0 48608 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_49_426
timestamp 1698431365
transform 1 0 49056 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_2
timestamp 1698431365
transform 1 0 1568 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_34
timestamp 1698431365
transform 1 0 5152 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_37
timestamp 1698431365
transform 1 0 5488 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_53
timestamp 1698431365
transform 1 0 7280 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_61
timestamp 1698431365
transform 1 0 8176 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_65
timestamp 1698431365
transform 1 0 8624 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_95
timestamp 1698431365
transform 1 0 11984 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_99
timestamp 1698431365
transform 1 0 12432 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_103
timestamp 1698431365
transform 1 0 12880 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_107
timestamp 1698431365
transform 1 0 13328 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_109
timestamp 1698431365
transform 1 0 13552 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_128
timestamp 1698431365
transform 1 0 15680 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_132
timestamp 1698431365
transform 1 0 16128 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_164
timestamp 1698431365
transform 1 0 19712 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_172
timestamp 1698431365
transform 1 0 20608 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_174
timestamp 1698431365
transform 1 0 20832 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_177
timestamp 1698431365
transform 1 0 21168 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_193
timestamp 1698431365
transform 1 0 22960 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_204
timestamp 1698431365
transform 1 0 24192 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_236
timestamp 1698431365
transform 1 0 27776 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_240
timestamp 1698431365
transform 1 0 28224 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_242
timestamp 1698431365
transform 1 0 28448 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_247
timestamp 1698431365
transform 1 0 29008 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_251
timestamp 1698431365
transform 1 0 29456 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_258
timestamp 1698431365
transform 1 0 30240 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_262
timestamp 1698431365
transform 1 0 30688 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_270
timestamp 1698431365
transform 1 0 31584 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_274
timestamp 1698431365
transform 1 0 32032 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_278
timestamp 1698431365
transform 1 0 32480 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_292
timestamp 1698431365
transform 1 0 34048 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_308
timestamp 1698431365
transform 1 0 35840 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_312
timestamp 1698431365
transform 1 0 36288 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_314
timestamp 1698431365
transform 1 0 36512 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_327
timestamp 1698431365
transform 1 0 37968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_329
timestamp 1698431365
transform 1 0 38192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_344
timestamp 1698431365
transform 1 0 39872 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_381
timestamp 1698431365
transform 1 0 44016 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_50_397
timestamp 1698431365
transform 1 0 45808 0 1 42336
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_50_429
timestamp 1698431365
transform 1 0 49392 0 1 42336
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_433
timestamp 1698431365
transform 1 0 49840 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_50_436
timestamp 1698431365
transform 1 0 50176 0 1 42336
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_50_452
timestamp 1698431365
transform 1 0 51968 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_50_454
timestamp 1698431365
transform 1 0 52192 0 1 42336
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_50_457
timestamp 1698431365
transform 1 0 52528 0 1 42336
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_51_2
timestamp 1698431365
transform 1 0 1568 0 -1 43904
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_66
timestamp 1698431365
transform 1 0 8736 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_72
timestamp 1698431365
transform 1 0 9408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_80
timestamp 1698431365
transform 1 0 10304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_103
timestamp 1698431365
transform 1 0 12880 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_111
timestamp 1698431365
transform 1 0 13776 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_120
timestamp 1698431365
transform 1 0 14784 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_136
timestamp 1698431365
transform 1 0 16576 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_142
timestamp 1698431365
transform 1 0 17248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_146
timestamp 1698431365
transform 1 0 17696 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_148
timestamp 1698431365
transform 1 0 17920 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_159
timestamp 1698431365
transform 1 0 19152 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_163
timestamp 1698431365
transform 1 0 19600 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_171
timestamp 1698431365
transform 1 0 20496 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_181
timestamp 1698431365
transform 1 0 21616 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_197
timestamp 1698431365
transform 1 0 23408 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_205
timestamp 1698431365
transform 1 0 24304 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_209
timestamp 1698431365
transform 1 0 24752 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_212
timestamp 1698431365
transform 1 0 25088 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_223
timestamp 1698431365
transform 1 0 26320 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_225
timestamp 1698431365
transform 1 0 26544 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_234
timestamp 1698431365
transform 1 0 27552 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_236
timestamp 1698431365
transform 1 0 27776 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_253
timestamp 1698431365
transform 1 0 29680 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_269
timestamp 1698431365
transform 1 0 31472 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_277
timestamp 1698431365
transform 1 0 32368 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_279
timestamp 1698431365
transform 1 0 32592 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_282
timestamp 1698431365
transform 1 0 32928 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_284
timestamp 1698431365
transform 1 0 33152 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_297
timestamp 1698431365
transform 1 0 34608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_301
timestamp 1698431365
transform 1 0 35056 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_338
timestamp 1698431365
transform 1 0 39200 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_346
timestamp 1698431365
transform 1 0 40096 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_51_352
timestamp 1698431365
transform 1 0 40768 0 -1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_51_384
timestamp 1698431365
transform 1 0 44352 0 -1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_51_392
timestamp 1698431365
transform 1 0 45248 0 -1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_396
timestamp 1698431365
transform 1 0 45696 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_51_402
timestamp 1698431365
transform 1 0 46368 0 -1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_422
timestamp 1698431365
transform 1 0 48608 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_424
timestamp 1698431365
transform 1 0 48832 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_51_433
timestamp 1698431365
transform 1 0 49840 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_51_435
timestamp 1698431365
transform 1 0 50064 0 -1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_2
timestamp 1698431365
transform 1 0 1568 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_34
timestamp 1698431365
transform 1 0 5152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_37
timestamp 1698431365
transform 1 0 5488 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_69
timestamp 1698431365
transform 1 0 9072 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_85
timestamp 1698431365
transform 1 0 10864 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_89
timestamp 1698431365
transform 1 0 11312 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_92
timestamp 1698431365
transform 1 0 11648 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_100
timestamp 1698431365
transform 1 0 12544 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_104
timestamp 1698431365
transform 1 0 12992 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_107
timestamp 1698431365
transform 1 0 13328 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_123
timestamp 1698431365
transform 1 0 15120 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_127
timestamp 1698431365
transform 1 0 15568 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_129
timestamp 1698431365
transform 1 0 15792 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_136
timestamp 1698431365
transform 1 0 16576 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_140
timestamp 1698431365
transform 1 0 17024 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_157
timestamp 1698431365
transform 1 0 18928 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_159
timestamp 1698431365
transform 1 0 19152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_172
timestamp 1698431365
transform 1 0 20608 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_174
timestamp 1698431365
transform 1 0 20832 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_177
timestamp 1698431365
transform 1 0 21168 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_181
timestamp 1698431365
transform 1 0 21616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_200
timestamp 1698431365
transform 1 0 23744 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_208
timestamp 1698431365
transform 1 0 24640 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_210
timestamp 1698431365
transform 1 0 24864 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_233
timestamp 1698431365
transform 1 0 27440 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_241
timestamp 1698431365
transform 1 0 28336 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_276
timestamp 1698431365
transform 1 0 32256 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_284
timestamp 1698431365
transform 1 0 33152 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_52_293
timestamp 1698431365
transform 1 0 34160 0 1 43904
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_317
timestamp 1698431365
transform 1 0 36848 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_335
timestamp 1698431365
transform 1 0 38864 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_52_367
timestamp 1698431365
transform 1 0 42448 0 1 43904
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_383
timestamp 1698431365
transform 1 0 44240 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_52_387
timestamp 1698431365
transform 1 0 44688 0 1 43904
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_431
timestamp 1698431365
transform 1 0 49616 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_433
timestamp 1698431365
transform 1 0 49840 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_436
timestamp 1698431365
transform 1 0 50176 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_444
timestamp 1698431365
transform 1 0 51072 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_52_452
timestamp 1698431365
transform 1 0 51968 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_52_454
timestamp 1698431365
transform 1 0 52192 0 1 43904
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_52_457
timestamp 1698431365
transform 1 0 52528 0 1 43904
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_53_2
timestamp 1698431365
transform 1 0 1568 0 -1 45472
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_66
timestamp 1698431365
transform 1 0 8736 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_72
timestamp 1698431365
transform 1 0 9408 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_80
timestamp 1698431365
transform 1 0 10304 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_84
timestamp 1698431365
transform 1 0 10752 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_86
timestamp 1698431365
transform 1 0 10976 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_101
timestamp 1698431365
transform 1 0 12656 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_109
timestamp 1698431365
transform 1 0 13552 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_111
timestamp 1698431365
transform 1 0 13776 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_122
timestamp 1698431365
transform 1 0 15008 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_124
timestamp 1698431365
transform 1 0 15232 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_127
timestamp 1698431365
transform 1 0 15568 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_135
timestamp 1698431365
transform 1 0 16464 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_139
timestamp 1698431365
transform 1 0 16912 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_142
timestamp 1698431365
transform 1 0 17248 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_146
timestamp 1698431365
transform 1 0 17696 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_161
timestamp 1698431365
transform 1 0 19376 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_53_165
timestamp 1698431365
transform 1 0 19824 0 -1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_181
timestamp 1698431365
transform 1 0 21616 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_185
timestamp 1698431365
transform 1 0 22064 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_187
timestamp 1698431365
transform 1 0 22288 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_200
timestamp 1698431365
transform 1 0 23744 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_204
timestamp 1698431365
transform 1 0 24192 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_206
timestamp 1698431365
transform 1 0 24416 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_209
timestamp 1698431365
transform 1 0 24752 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_212
timestamp 1698431365
transform 1 0 25088 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_216
timestamp 1698431365
transform 1 0 25536 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_218
timestamp 1698431365
transform 1 0 25760 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_53_223
timestamp 1698431365
transform 1 0 26320 0 -1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_255
timestamp 1698431365
transform 1 0 29904 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_53_263
timestamp 1698431365
transform 1 0 30800 0 -1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_267
timestamp 1698431365
transform 1 0 31248 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_278
timestamp 1698431365
transform 1 0 32480 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_282
timestamp 1698431365
transform 1 0 32928 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_316
timestamp 1698431365
transform 1 0 36736 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_342
timestamp 1698431365
transform 1 0 39648 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_53_361
timestamp 1698431365
transform 1 0 41776 0 -1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_369
timestamp 1698431365
transform 1 0 42672 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_53_376
timestamp 1698431365
transform 1 0 43456 0 -1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_406
timestamp 1698431365
transform 1 0 46816 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_410
timestamp 1698431365
transform 1 0 47264 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_53_437
timestamp 1698431365
transform 1 0 50288 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_2
timestamp 1698431365
transform 1 0 1568 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_34
timestamp 1698431365
transform 1 0 5152 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_37
timestamp 1698431365
transform 1 0 5488 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_53
timestamp 1698431365
transform 1 0 7280 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_61
timestamp 1698431365
transform 1 0 8176 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_63
timestamp 1698431365
transform 1 0 8400 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_93
timestamp 1698431365
transform 1 0 11760 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_102
timestamp 1698431365
transform 1 0 12768 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_104
timestamp 1698431365
transform 1 0 12992 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_107
timestamp 1698431365
transform 1 0 13328 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_111
timestamp 1698431365
transform 1 0 13776 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_125
timestamp 1698431365
transform 1 0 15344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_127
timestamp 1698431365
transform 1 0 15568 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_157
timestamp 1698431365
transform 1 0 18928 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_161
timestamp 1698431365
transform 1 0 19376 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_169
timestamp 1698431365
transform 1 0 20272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_173
timestamp 1698431365
transform 1 0 20720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_177
timestamp 1698431365
transform 1 0 21168 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_195
timestamp 1698431365
transform 1 0 23184 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_199
timestamp 1698431365
transform 1 0 23632 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_213
timestamp 1698431365
transform 1 0 25200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_217
timestamp 1698431365
transform 1 0 25648 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_233
timestamp 1698431365
transform 1 0 27440 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_241
timestamp 1698431365
transform 1 0 28336 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_247
timestamp 1698431365
transform 1 0 29008 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_279
timestamp 1698431365
transform 1 0 32592 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_287
timestamp 1698431365
transform 1 0 33488 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_289
timestamp 1698431365
transform 1 0 33712 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_296
timestamp 1698431365
transform 1 0 34496 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_312
timestamp 1698431365
transform 1 0 36288 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_314
timestamp 1698431365
transform 1 0 36512 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_330
timestamp 1698431365
transform 1 0 38304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_334
timestamp 1698431365
transform 1 0 38752 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_338
timestamp 1698431365
transform 1 0 39200 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_352
timestamp 1698431365
transform 1 0 40768 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_54_384
timestamp 1698431365
transform 1 0 44352 0 1 45472
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_54_387
timestamp 1698431365
transform 1 0 44688 0 1 45472
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_54_419
timestamp 1698431365
transform 1 0 48272 0 1 45472
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_423
timestamp 1698431365
transform 1 0 48720 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_54_429
timestamp 1698431365
transform 1 0 49392 0 1 45472
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_445
timestamp 1698431365
transform 1 0 51184 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_54_453
timestamp 1698431365
transform 1 0 52080 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_54_457
timestamp 1698431365
transform 1 0 52528 0 1 45472
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_55_2
timestamp 1698431365
transform 1 0 1568 0 -1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_66
timestamp 1698431365
transform 1 0 8736 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_72
timestamp 1698431365
transform 1 0 9408 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_88
timestamp 1698431365
transform 1 0 11200 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_92
timestamp 1698431365
transform 1 0 11648 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_100
timestamp 1698431365
transform 1 0 12544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_125
timestamp 1698431365
transform 1 0 15344 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_133
timestamp 1698431365
transform 1 0 16240 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_137
timestamp 1698431365
transform 1 0 16688 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_139
timestamp 1698431365
transform 1 0 16912 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_142
timestamp 1698431365
transform 1 0 17248 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_150
timestamp 1698431365
transform 1 0 18144 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_154
timestamp 1698431365
transform 1 0 18592 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_171
timestamp 1698431365
transform 1 0 20496 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_212
timestamp 1698431365
transform 1 0 25088 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_228
timestamp 1698431365
transform 1 0 26880 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_230
timestamp 1698431365
transform 1 0 27104 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_236
timestamp 1698431365
transform 1 0 27776 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_252
timestamp 1698431365
transform 1 0 29568 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_254
timestamp 1698431365
transform 1 0 29792 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_268
timestamp 1698431365
transform 1 0 31360 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_278
timestamp 1698431365
transform 1 0 32480 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_282
timestamp 1698431365
transform 1 0 32928 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_292
timestamp 1698431365
transform 1 0 34048 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_300
timestamp 1698431365
transform 1 0 34944 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_302
timestamp 1698431365
transform 1 0 35168 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_340
timestamp 1698431365
transform 1 0 39424 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_55_352
timestamp 1698431365
transform 1 0 40768 0 -1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_55_368
timestamp 1698431365
transform 1 0 42560 0 -1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_376
timestamp 1698431365
transform 1 0 43456 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_380
timestamp 1698431365
transform 1 0 43904 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_55_382
timestamp 1698431365
transform 1 0 44128 0 -1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_412
timestamp 1698431365
transform 1 0 47488 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_55_416
timestamp 1698431365
transform 1 0 47936 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_55_430
timestamp 1698431365
transform 1 0 49504 0 -1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_2
timestamp 1698431365
transform 1 0 1568 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_34
timestamp 1698431365
transform 1 0 5152 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_56_37
timestamp 1698431365
transform 1 0 5488 0 1 47040
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_101
timestamp 1698431365
transform 1 0 12656 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_107
timestamp 1698431365
transform 1 0 13328 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_56_119
timestamp 1698431365
transform 1 0 14672 0 1 47040
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_151
timestamp 1698431365
transform 1 0 18256 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_165
timestamp 1698431365
transform 1 0 19824 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_173
timestamp 1698431365
transform 1 0 20720 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_177
timestamp 1698431365
transform 1 0 21168 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_193
timestamp 1698431365
transform 1 0 22960 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_197
timestamp 1698431365
transform 1 0 23408 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_242
timestamp 1698431365
transform 1 0 28448 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_244
timestamp 1698431365
transform 1 0 28672 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_305
timestamp 1698431365
transform 1 0 35504 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_309
timestamp 1698431365
transform 1 0 35952 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_313
timestamp 1698431365
transform 1 0 36400 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_317
timestamp 1698431365
transform 1 0 36848 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_325
timestamp 1698431365
transform 1 0 37744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_329
timestamp 1698431365
transform 1 0 38192 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_331
timestamp 1698431365
transform 1 0 38416 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_334
timestamp 1698431365
transform 1 0 38752 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_350
timestamp 1698431365
transform 1 0 40544 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_367
timestamp 1698431365
transform 1 0 42448 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_374
timestamp 1698431365
transform 1 0 43232 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_382
timestamp 1698431365
transform 1 0 44128 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_384
timestamp 1698431365
transform 1 0 44352 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_387
timestamp 1698431365
transform 1 0 44688 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_395
timestamp 1698431365
transform 1 0 45584 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_399
timestamp 1698431365
transform 1 0 46032 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_56_402
timestamp 1698431365
transform 1 0 46368 0 1 47040
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_418
timestamp 1698431365
transform 1 0 48160 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_56_446
timestamp 1698431365
transform 1 0 51296 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_56_450
timestamp 1698431365
transform 1 0 51744 0 1 47040
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_56_454
timestamp 1698431365
transform 1 0 52192 0 1 47040
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_56_457
timestamp 1698431365
transform 1 0 52528 0 1 47040
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_2
timestamp 1698431365
transform 1 0 1568 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_66
timestamp 1698431365
transform 1 0 8736 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_57_72
timestamp 1698431365
transform 1 0 9408 0 -1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_136
timestamp 1698431365
transform 1 0 16576 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_142
timestamp 1698431365
transform 1 0 17248 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_158
timestamp 1698431365
transform 1 0 19040 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_160
timestamp 1698431365
transform 1 0 19264 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_192
timestamp 1698431365
transform 1 0 22848 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_196
timestamp 1698431365
transform 1 0 23296 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_200
timestamp 1698431365
transform 1 0 23744 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_209
timestamp 1698431365
transform 1 0 24752 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_220
timestamp 1698431365
transform 1 0 25984 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_232
timestamp 1698431365
transform 1 0 27328 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_236
timestamp 1698431365
transform 1 0 27776 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_268
timestamp 1698431365
transform 1 0 31360 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_275
timestamp 1698431365
transform 1 0 32144 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_279
timestamp 1698431365
transform 1 0 32592 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_57_282
timestamp 1698431365
transform 1 0 32928 0 -1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_57_314
timestamp 1698431365
transform 1 0 36512 0 -1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_330
timestamp 1698431365
transform 1 0 38304 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_338
timestamp 1698431365
transform 1 0 39200 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_348
timestamp 1698431365
transform 1 0 40320 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_352
timestamp 1698431365
transform 1 0 40768 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_57_356
timestamp 1698431365
transform 1 0 41216 0 -1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_57_360
timestamp 1698431365
transform 1 0 41664 0 -1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_398
timestamp 1698431365
transform 1 0 45920 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_57_410
timestamp 1698431365
transform 1 0 47264 0 -1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_430
timestamp 1698431365
transform 1 0 49504 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_57_437
timestamp 1698431365
transform 1 0 50288 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_2
timestamp 1698431365
transform 1 0 1568 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_34
timestamp 1698431365
transform 1 0 5152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_58_37
timestamp 1698431365
transform 1 0 5488 0 1 48608
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_101
timestamp 1698431365
transform 1 0 12656 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_136
timestamp 1698431365
transform 1 0 16576 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_140
timestamp 1698431365
transform 1 0 17024 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_148
timestamp 1698431365
transform 1 0 17920 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_155
timestamp 1698431365
transform 1 0 18704 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_159
timestamp 1698431365
transform 1 0 19152 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_171
timestamp 1698431365
transform 1 0 20496 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_177
timestamp 1698431365
transform 1 0 21168 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_209
timestamp 1698431365
transform 1 0 24752 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_225
timestamp 1698431365
transform 1 0 26544 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_233
timestamp 1698431365
transform 1 0 27440 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_241
timestamp 1698431365
transform 1 0 28336 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_247
timestamp 1698431365
transform 1 0 29008 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_263
timestamp 1698431365
transform 1 0 30800 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_58_266
timestamp 1698431365
transform 1 0 31136 0 1 48608
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_298
timestamp 1698431365
transform 1 0 34720 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_306
timestamp 1698431365
transform 1 0 35616 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_314
timestamp 1698431365
transform 1 0 36512 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_317
timestamp 1698431365
transform 1 0 36848 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_321
timestamp 1698431365
transform 1 0 37296 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_325
timestamp 1698431365
transform 1 0 37744 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_335
timestamp 1698431365
transform 1 0 38864 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_351
timestamp 1698431365
transform 1 0 40656 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_58_361
timestamp 1698431365
transform 1 0 41776 0 1 48608
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_377
timestamp 1698431365
transform 1 0 43568 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_387
timestamp 1698431365
transform 1 0 44688 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_58_395
timestamp 1698431365
transform 1 0 45584 0 1 48608
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_58_399
timestamp 1698431365
transform 1 0 46032 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_58_401
timestamp 1698431365
transform 1 0 46256 0 1 48608
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_411
timestamp 1698431365
transform 1 0 47376 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_58_457
timestamp 1698431365
transform 1 0 52528 0 1 48608
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_2
timestamp 1698431365
transform 1 0 1568 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_66
timestamp 1698431365
transform 1 0 8736 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_59_72
timestamp 1698431365
transform 1 0 9408 0 -1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_136
timestamp 1698431365
transform 1 0 16576 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_150
timestamp 1698431365
transform 1 0 18144 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_158
timestamp 1698431365
transform 1 0 19040 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_162
timestamp 1698431365
transform 1 0 19488 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_204
timestamp 1698431365
transform 1 0 24192 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_208
timestamp 1698431365
transform 1 0 24640 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_221
timestamp 1698431365
transform 1 0 26096 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_276
timestamp 1698431365
transform 1 0 32256 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_282
timestamp 1698431365
transform 1 0 32928 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_319
timestamp 1698431365
transform 1 0 37072 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_335
timestamp 1698431365
transform 1 0 38864 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_343
timestamp 1698431365
transform 1 0 39760 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_347
timestamp 1698431365
transform 1 0 40208 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_59_349
timestamp 1698431365
transform 1 0 40432 0 -1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_59_352
timestamp 1698431365
transform 1 0 40768 0 -1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_59_366
timestamp 1698431365
transform 1 0 42336 0 -1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_59_398
timestamp 1698431365
transform 1 0 45920 0 -1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_59_414
timestamp 1698431365
transform 1 0 47712 0 -1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_59_432
timestamp 1698431365
transform 1 0 49728 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_60_2
timestamp 1698431365
transform 1 0 1568 0 1 50176
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_34
timestamp 1698431365
transform 1 0 5152 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_60_37
timestamp 1698431365
transform 1 0 5488 0 1 50176
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_101
timestamp 1698431365
transform 1 0 12656 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_107
timestamp 1698431365
transform 1 0 13328 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_123
timestamp 1698431365
transform 1 0 15120 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_125
timestamp 1698431365
transform 1 0 15344 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_155
timestamp 1698431365
transform 1 0 18704 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_159
timestamp 1698431365
transform 1 0 19152 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_177
timestamp 1698431365
transform 1 0 21168 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_193
timestamp 1698431365
transform 1 0 22960 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_214
timestamp 1698431365
transform 1 0 25312 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_238
timestamp 1698431365
transform 1 0 28000 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_242
timestamp 1698431365
transform 1 0 28448 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_244
timestamp 1698431365
transform 1 0 28672 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_247
timestamp 1698431365
transform 1 0 29008 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_263
timestamp 1698431365
transform 1 0 30800 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_293
timestamp 1698431365
transform 1 0 34160 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_60_297
timestamp 1698431365
transform 1 0 34608 0 1 50176
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_313
timestamp 1698431365
transform 1 0 36400 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_317
timestamp 1698431365
transform 1 0 36848 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_350
timestamp 1698431365
transform 1 0 40544 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_354
timestamp 1698431365
transform 1 0 40992 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_384
timestamp 1698431365
transform 1 0 44352 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_387
timestamp 1698431365
transform 1 0 44688 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_60_391
timestamp 1698431365
transform 1 0 45136 0 1 50176
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_60_421
timestamp 1698431365
transform 1 0 48496 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_60_425
timestamp 1698431365
transform 1 0 48944 0 1 50176
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_60_457
timestamp 1698431365
transform 1 0 52528 0 1 50176
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_2
timestamp 1698431365
transform 1 0 1568 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_36
timestamp 1698431365
transform 1 0 5376 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_70
timestamp 1698431365
transform 1 0 9184 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_104
timestamp 1698431365
transform 1 0 12992 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_138
timestamp 1698431365
transform 1 0 16800 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_172
timestamp 1698431365
transform 1 0 20608 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_206
timestamp 1698431365
transform 1 0 24416 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_240
timestamp 1698431365
transform 1 0 28224 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_274
timestamp 1698431365
transform 1 0 32032 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_308
timestamp 1698431365
transform 1 0 35840 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_342
timestamp 1698431365
transform 1 0 39648 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_350
timestamp 1698431365
transform 1 0 40544 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_354
timestamp 1698431365
transform 1 0 40992 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_363
timestamp 1698431365
transform 1 0 42000 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_371
timestamp 1698431365
transform 1 0 42896 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_373
timestamp 1698431365
transform 1 0 43120 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_61_376
timestamp 1698431365
transform 1 0 43456 0 -1 51744
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_61_410
timestamp 1698431365
transform 1 0 47264 0 -1 51744
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_426
timestamp 1698431365
transform 1 0 49056 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_61_430
timestamp 1698431365
transform 1 0 49504 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_61_452
timestamp 1698431365
transform 1 0 51968 0 -1 51744
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_61_460
timestamp 1698431365
transform 1 0 52864 0 -1 51744
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_61_464
timestamp 1698431365
transform 1 0 53312 0 -1 51744
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input1
timestamp 1698431365
transform 1 0 39648 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input2
timestamp 1698431365
transform -1 0 53424 0 1 3136
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input3
timestamp 1698431365
transform -1 0 52304 0 1 6272
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input4
timestamp 1698431365
transform -1 0 53424 0 -1 9408
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input5
timestamp 1698431365
transform 1 0 43456 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input6
timestamp 1698431365
transform -1 0 47936 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input7
timestamp 1698431365
transform -1 0 53424 0 1 10976
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  input8
timestamp 1698431365
transform -1 0 53424 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input9
timestamp 1698431365
transform -1 0 53424 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input10
timestamp 1698431365
transform -1 0 53424 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input11
timestamp 1698431365
transform -1 0 53424 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input12
timestamp 1698431365
transform -1 0 53424 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input13
timestamp 1698431365
transform -1 0 53424 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input14
timestamp 1698431365
transform -1 0 53424 0 1 29792
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  input15
timestamp 1698431365
transform 1 0 2800 0 1 3136
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  input16
timestamp 1698431365
transform 1 0 41328 0 -1 51744
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 35840 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698431365
transform 1 0 50512 0 -1 32928
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698431365
transform 1 0 50512 0 -1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698431365
transform 1 0 50512 0 -1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698431365
transform 1 0 49392 0 1 40768
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698431365
transform 1 0 50512 0 -1 45472
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698431365
transform 1 0 50512 0 -1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698431365
transform 1 0 49392 0 1 48608
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698431365
transform -1 0 52304 0 1 50176
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698431365
transform -1 0 12096 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output27
timestamp 1698431365
transform -1 0 14672 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output28
timestamp 1698431365
transform 1 0 47936 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_62 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698431365
transform -1 0 53648 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_63
timestamp 1698431365
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698431365
transform -1 0 53648 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_64
timestamp 1698431365
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698431365
transform -1 0 53648 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_65
timestamp 1698431365
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698431365
transform -1 0 53648 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_66
timestamp 1698431365
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698431365
transform -1 0 53648 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_67
timestamp 1698431365
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698431365
transform -1 0 53648 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_68
timestamp 1698431365
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698431365
transform -1 0 53648 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_69
timestamp 1698431365
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698431365
transform -1 0 53648 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_70
timestamp 1698431365
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698431365
transform -1 0 53648 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_71
timestamp 1698431365
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698431365
transform -1 0 53648 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_72
timestamp 1698431365
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698431365
transform -1 0 53648 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_73
timestamp 1698431365
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698431365
transform -1 0 53648 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_74
timestamp 1698431365
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698431365
transform -1 0 53648 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_75
timestamp 1698431365
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698431365
transform -1 0 53648 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_76
timestamp 1698431365
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698431365
transform -1 0 53648 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_77
timestamp 1698431365
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698431365
transform -1 0 53648 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_78
timestamp 1698431365
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698431365
transform -1 0 53648 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_79
timestamp 1698431365
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698431365
transform -1 0 53648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_80
timestamp 1698431365
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698431365
transform -1 0 53648 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_81
timestamp 1698431365
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698431365
transform -1 0 53648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_82
timestamp 1698431365
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698431365
transform -1 0 53648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_83
timestamp 1698431365
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698431365
transform -1 0 53648 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_84
timestamp 1698431365
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698431365
transform -1 0 53648 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_85
timestamp 1698431365
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698431365
transform -1 0 53648 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_86
timestamp 1698431365
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698431365
transform -1 0 53648 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_87
timestamp 1698431365
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698431365
transform -1 0 53648 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_88
timestamp 1698431365
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698431365
transform -1 0 53648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_89
timestamp 1698431365
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698431365
transform -1 0 53648 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_90
timestamp 1698431365
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698431365
transform -1 0 53648 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_91
timestamp 1698431365
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698431365
transform -1 0 53648 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_92
timestamp 1698431365
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698431365
transform -1 0 53648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_93
timestamp 1698431365
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698431365
transform -1 0 53648 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_94
timestamp 1698431365
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698431365
transform -1 0 53648 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_95
timestamp 1698431365
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698431365
transform -1 0 53648 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_96
timestamp 1698431365
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698431365
transform -1 0 53648 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_97
timestamp 1698431365
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698431365
transform -1 0 53648 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_98
timestamp 1698431365
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698431365
transform -1 0 53648 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_99
timestamp 1698431365
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698431365
transform -1 0 53648 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_100
timestamp 1698431365
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698431365
transform -1 0 53648 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_101
timestamp 1698431365
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698431365
transform -1 0 53648 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_102
timestamp 1698431365
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698431365
transform -1 0 53648 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_103
timestamp 1698431365
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698431365
transform -1 0 53648 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_104
timestamp 1698431365
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698431365
transform -1 0 53648 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_105
timestamp 1698431365
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698431365
transform -1 0 53648 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_106
timestamp 1698431365
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698431365
transform -1 0 53648 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Left_107
timestamp 1698431365
transform 1 0 1344 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_45_Right_45
timestamp 1698431365
transform -1 0 53648 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Left_108
timestamp 1698431365
transform 1 0 1344 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_46_Right_46
timestamp 1698431365
transform -1 0 53648 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Left_109
timestamp 1698431365
transform 1 0 1344 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_47_Right_47
timestamp 1698431365
transform -1 0 53648 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Left_110
timestamp 1698431365
transform 1 0 1344 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_48_Right_48
timestamp 1698431365
transform -1 0 53648 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Left_111
timestamp 1698431365
transform 1 0 1344 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_49_Right_49
timestamp 1698431365
transform -1 0 53648 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Left_112
timestamp 1698431365
transform 1 0 1344 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_50_Right_50
timestamp 1698431365
transform -1 0 53648 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Left_113
timestamp 1698431365
transform 1 0 1344 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_51_Right_51
timestamp 1698431365
transform -1 0 53648 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Left_114
timestamp 1698431365
transform 1 0 1344 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_52_Right_52
timestamp 1698431365
transform -1 0 53648 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Left_115
timestamp 1698431365
transform 1 0 1344 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_53_Right_53
timestamp 1698431365
transform -1 0 53648 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Left_116
timestamp 1698431365
transform 1 0 1344 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_54_Right_54
timestamp 1698431365
transform -1 0 53648 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Left_117
timestamp 1698431365
transform 1 0 1344 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_55_Right_55
timestamp 1698431365
transform -1 0 53648 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Left_118
timestamp 1698431365
transform 1 0 1344 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_56_Right_56
timestamp 1698431365
transform -1 0 53648 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Left_119
timestamp 1698431365
transform 1 0 1344 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_57_Right_57
timestamp 1698431365
transform -1 0 53648 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Left_120
timestamp 1698431365
transform 1 0 1344 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_58_Right_58
timestamp 1698431365
transform -1 0 53648 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Left_121
timestamp 1698431365
transform 1 0 1344 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_59_Right_59
timestamp 1698431365
transform -1 0 53648 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Left_122
timestamp 1698431365
transform 1 0 1344 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_60_Right_60
timestamp 1698431365
transform -1 0 53648 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Left_123
timestamp 1698431365
transform 1 0 1344 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_61_Right_61
timestamp 1698431365
transform -1 0 53648 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_29 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 21168 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_30
timestamp 1698431365
transform -1 0 25648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  serial_ports_31
timestamp 1698431365
transform -1 0 17248 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  serial_ports_32 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform -1 0 30128 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_124 $PDKPATH/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698431365
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_125
timestamp 1698431365
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_126
timestamp 1698431365
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_127
timestamp 1698431365
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_128
timestamp 1698431365
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_129
timestamp 1698431365
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_130
timestamp 1698431365
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_131
timestamp 1698431365
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_132
timestamp 1698431365
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_133
timestamp 1698431365
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_134
timestamp 1698431365
transform 1 0 43232 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_135
timestamp 1698431365
transform 1 0 47040 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_136
timestamp 1698431365
transform 1 0 50848 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_137
timestamp 1698431365
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_138
timestamp 1698431365
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_139
timestamp 1698431365
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_140
timestamp 1698431365
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_141
timestamp 1698431365
transform 1 0 40544 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_142
timestamp 1698431365
transform 1 0 48384 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_143
timestamp 1698431365
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_144
timestamp 1698431365
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_145
timestamp 1698431365
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_146
timestamp 1698431365
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_147
timestamp 1698431365
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_148
timestamp 1698431365
transform 1 0 44464 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_149
timestamp 1698431365
transform 1 0 52304 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_150
timestamp 1698431365
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_151
timestamp 1698431365
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_152
timestamp 1698431365
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_153
timestamp 1698431365
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_154
timestamp 1698431365
transform 1 0 40544 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_155
timestamp 1698431365
transform 1 0 48384 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_156
timestamp 1698431365
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_157
timestamp 1698431365
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_158
timestamp 1698431365
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_159
timestamp 1698431365
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_160
timestamp 1698431365
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_161
timestamp 1698431365
transform 1 0 44464 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_162
timestamp 1698431365
transform 1 0 52304 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_163
timestamp 1698431365
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_164
timestamp 1698431365
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_165
timestamp 1698431365
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_166
timestamp 1698431365
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_167
timestamp 1698431365
transform 1 0 40544 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_168
timestamp 1698431365
transform 1 0 48384 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_169
timestamp 1698431365
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_170
timestamp 1698431365
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_171
timestamp 1698431365
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_172
timestamp 1698431365
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_173
timestamp 1698431365
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_174
timestamp 1698431365
transform 1 0 44464 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_175
timestamp 1698431365
transform 1 0 52304 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_176
timestamp 1698431365
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_177
timestamp 1698431365
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_178
timestamp 1698431365
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_179
timestamp 1698431365
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_180
timestamp 1698431365
transform 1 0 40544 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_181
timestamp 1698431365
transform 1 0 48384 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_182
timestamp 1698431365
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_183
timestamp 1698431365
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_184
timestamp 1698431365
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_185
timestamp 1698431365
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_186
timestamp 1698431365
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_187
timestamp 1698431365
transform 1 0 44464 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_188
timestamp 1698431365
transform 1 0 52304 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_189
timestamp 1698431365
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_190
timestamp 1698431365
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_191
timestamp 1698431365
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_192
timestamp 1698431365
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_193
timestamp 1698431365
transform 1 0 40544 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_194
timestamp 1698431365
transform 1 0 48384 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_195
timestamp 1698431365
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_196
timestamp 1698431365
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_197
timestamp 1698431365
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_198
timestamp 1698431365
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_199
timestamp 1698431365
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_200
timestamp 1698431365
transform 1 0 44464 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_201
timestamp 1698431365
transform 1 0 52304 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_202
timestamp 1698431365
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_203
timestamp 1698431365
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_204
timestamp 1698431365
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_205
timestamp 1698431365
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_206
timestamp 1698431365
transform 1 0 40544 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_207
timestamp 1698431365
transform 1 0 48384 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_208
timestamp 1698431365
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_209
timestamp 1698431365
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_210
timestamp 1698431365
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_211
timestamp 1698431365
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_212
timestamp 1698431365
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_213
timestamp 1698431365
transform 1 0 44464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_214
timestamp 1698431365
transform 1 0 52304 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_215
timestamp 1698431365
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_216
timestamp 1698431365
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_217
timestamp 1698431365
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_218
timestamp 1698431365
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_219
timestamp 1698431365
transform 1 0 40544 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_220
timestamp 1698431365
transform 1 0 48384 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_221
timestamp 1698431365
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_222
timestamp 1698431365
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_223
timestamp 1698431365
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_224
timestamp 1698431365
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_225
timestamp 1698431365
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_226
timestamp 1698431365
transform 1 0 44464 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_227
timestamp 1698431365
transform 1 0 52304 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_228
timestamp 1698431365
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_229
timestamp 1698431365
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_230
timestamp 1698431365
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_231
timestamp 1698431365
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_232
timestamp 1698431365
transform 1 0 40544 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_233
timestamp 1698431365
transform 1 0 48384 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_234
timestamp 1698431365
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_235
timestamp 1698431365
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_236
timestamp 1698431365
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_237
timestamp 1698431365
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_238
timestamp 1698431365
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_239
timestamp 1698431365
transform 1 0 44464 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_240
timestamp 1698431365
transform 1 0 52304 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_241
timestamp 1698431365
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_242
timestamp 1698431365
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_243
timestamp 1698431365
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_244
timestamp 1698431365
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_245
timestamp 1698431365
transform 1 0 40544 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_246
timestamp 1698431365
transform 1 0 48384 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_247
timestamp 1698431365
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_248
timestamp 1698431365
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_249
timestamp 1698431365
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_250
timestamp 1698431365
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_251
timestamp 1698431365
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_252
timestamp 1698431365
transform 1 0 44464 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_253
timestamp 1698431365
transform 1 0 52304 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_254
timestamp 1698431365
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_255
timestamp 1698431365
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_256
timestamp 1698431365
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_257
timestamp 1698431365
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_258
timestamp 1698431365
transform 1 0 40544 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_259
timestamp 1698431365
transform 1 0 48384 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_260
timestamp 1698431365
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_261
timestamp 1698431365
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_262
timestamp 1698431365
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_263
timestamp 1698431365
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_264
timestamp 1698431365
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_265
timestamp 1698431365
transform 1 0 44464 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_266
timestamp 1698431365
transform 1 0 52304 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_267
timestamp 1698431365
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_268
timestamp 1698431365
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_269
timestamp 1698431365
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_270
timestamp 1698431365
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_271
timestamp 1698431365
transform 1 0 40544 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_272
timestamp 1698431365
transform 1 0 48384 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_273
timestamp 1698431365
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_274
timestamp 1698431365
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_275
timestamp 1698431365
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_276
timestamp 1698431365
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_277
timestamp 1698431365
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_278
timestamp 1698431365
transform 1 0 44464 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_279
timestamp 1698431365
transform 1 0 52304 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_280
timestamp 1698431365
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_281
timestamp 1698431365
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_282
timestamp 1698431365
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_283
timestamp 1698431365
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_284
timestamp 1698431365
transform 1 0 40544 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_285
timestamp 1698431365
transform 1 0 48384 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_286
timestamp 1698431365
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_287
timestamp 1698431365
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_288
timestamp 1698431365
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_289
timestamp 1698431365
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_290
timestamp 1698431365
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_291
timestamp 1698431365
transform 1 0 44464 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_292
timestamp 1698431365
transform 1 0 52304 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_293
timestamp 1698431365
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_294
timestamp 1698431365
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_295
timestamp 1698431365
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_296
timestamp 1698431365
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_297
timestamp 1698431365
transform 1 0 40544 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_298
timestamp 1698431365
transform 1 0 48384 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_299
timestamp 1698431365
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_300
timestamp 1698431365
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_301
timestamp 1698431365
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_302
timestamp 1698431365
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_303
timestamp 1698431365
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_304
timestamp 1698431365
transform 1 0 44464 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_305
timestamp 1698431365
transform 1 0 52304 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_306
timestamp 1698431365
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_307
timestamp 1698431365
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_308
timestamp 1698431365
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_309
timestamp 1698431365
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_310
timestamp 1698431365
transform 1 0 40544 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_311
timestamp 1698431365
transform 1 0 48384 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_312
timestamp 1698431365
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_313
timestamp 1698431365
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_314
timestamp 1698431365
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_315
timestamp 1698431365
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_316
timestamp 1698431365
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_317
timestamp 1698431365
transform 1 0 44464 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_318
timestamp 1698431365
transform 1 0 52304 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_319
timestamp 1698431365
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_320
timestamp 1698431365
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_321
timestamp 1698431365
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_322
timestamp 1698431365
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_323
timestamp 1698431365
transform 1 0 40544 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_324
timestamp 1698431365
transform 1 0 48384 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_325
timestamp 1698431365
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_326
timestamp 1698431365
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_327
timestamp 1698431365
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_328
timestamp 1698431365
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_329
timestamp 1698431365
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_330
timestamp 1698431365
transform 1 0 44464 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_331
timestamp 1698431365
transform 1 0 52304 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_332
timestamp 1698431365
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_333
timestamp 1698431365
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_334
timestamp 1698431365
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_335
timestamp 1698431365
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_336
timestamp 1698431365
transform 1 0 40544 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_337
timestamp 1698431365
transform 1 0 48384 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_338
timestamp 1698431365
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_339
timestamp 1698431365
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_340
timestamp 1698431365
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_341
timestamp 1698431365
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_342
timestamp 1698431365
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_343
timestamp 1698431365
transform 1 0 44464 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_344
timestamp 1698431365
transform 1 0 52304 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_345
timestamp 1698431365
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_346
timestamp 1698431365
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_347
timestamp 1698431365
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_348
timestamp 1698431365
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_349
timestamp 1698431365
transform 1 0 40544 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_350
timestamp 1698431365
transform 1 0 48384 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_351
timestamp 1698431365
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_352
timestamp 1698431365
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_353
timestamp 1698431365
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_354
timestamp 1698431365
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_355
timestamp 1698431365
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_356
timestamp 1698431365
transform 1 0 44464 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_357
timestamp 1698431365
transform 1 0 52304 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_358
timestamp 1698431365
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_359
timestamp 1698431365
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_360
timestamp 1698431365
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_361
timestamp 1698431365
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_362
timestamp 1698431365
transform 1 0 40544 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_363
timestamp 1698431365
transform 1 0 48384 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_364
timestamp 1698431365
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_365
timestamp 1698431365
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_366
timestamp 1698431365
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_367
timestamp 1698431365
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_368
timestamp 1698431365
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_369
timestamp 1698431365
transform 1 0 44464 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_370
timestamp 1698431365
transform 1 0 52304 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_371
timestamp 1698431365
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_372
timestamp 1698431365
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_373
timestamp 1698431365
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_374
timestamp 1698431365
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_375
timestamp 1698431365
transform 1 0 40544 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_376
timestamp 1698431365
transform 1 0 48384 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_377
timestamp 1698431365
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_378
timestamp 1698431365
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_379
timestamp 1698431365
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_380
timestamp 1698431365
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_381
timestamp 1698431365
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_382
timestamp 1698431365
transform 1 0 44464 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_383
timestamp 1698431365
transform 1 0 52304 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_384
timestamp 1698431365
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_385
timestamp 1698431365
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_386
timestamp 1698431365
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_387
timestamp 1698431365
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_388
timestamp 1698431365
transform 1 0 40544 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_389
timestamp 1698431365
transform 1 0 48384 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_390
timestamp 1698431365
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_391
timestamp 1698431365
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_392
timestamp 1698431365
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_393
timestamp 1698431365
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_394
timestamp 1698431365
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_395
timestamp 1698431365
transform 1 0 44464 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_396
timestamp 1698431365
transform 1 0 52304 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_397
timestamp 1698431365
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_398
timestamp 1698431365
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_399
timestamp 1698431365
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_400
timestamp 1698431365
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_401
timestamp 1698431365
transform 1 0 40544 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_402
timestamp 1698431365
transform 1 0 48384 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_403
timestamp 1698431365
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_404
timestamp 1698431365
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_405
timestamp 1698431365
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_406
timestamp 1698431365
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_407
timestamp 1698431365
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_408
timestamp 1698431365
transform 1 0 44464 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_409
timestamp 1698431365
transform 1 0 52304 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_410
timestamp 1698431365
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_411
timestamp 1698431365
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_412
timestamp 1698431365
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_413
timestamp 1698431365
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_414
timestamp 1698431365
transform 1 0 40544 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_415
timestamp 1698431365
transform 1 0 48384 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_416
timestamp 1698431365
transform 1 0 5264 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_417
timestamp 1698431365
transform 1 0 13104 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_418
timestamp 1698431365
transform 1 0 20944 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_419
timestamp 1698431365
transform 1 0 28784 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_420
timestamp 1698431365
transform 1 0 36624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_421
timestamp 1698431365
transform 1 0 44464 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_422
timestamp 1698431365
transform 1 0 52304 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_423
timestamp 1698431365
transform 1 0 9184 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_424
timestamp 1698431365
transform 1 0 17024 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_425
timestamp 1698431365
transform 1 0 24864 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_426
timestamp 1698431365
transform 1 0 32704 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_427
timestamp 1698431365
transform 1 0 40544 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_45_428
timestamp 1698431365
transform 1 0 48384 0 -1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_429
timestamp 1698431365
transform 1 0 5264 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_430
timestamp 1698431365
transform 1 0 13104 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_431
timestamp 1698431365
transform 1 0 20944 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_432
timestamp 1698431365
transform 1 0 28784 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_433
timestamp 1698431365
transform 1 0 36624 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_434
timestamp 1698431365
transform 1 0 44464 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_46_435
timestamp 1698431365
transform 1 0 52304 0 1 39200
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_436
timestamp 1698431365
transform 1 0 9184 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_437
timestamp 1698431365
transform 1 0 17024 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_438
timestamp 1698431365
transform 1 0 24864 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_439
timestamp 1698431365
transform 1 0 32704 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_440
timestamp 1698431365
transform 1 0 40544 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_47_441
timestamp 1698431365
transform 1 0 48384 0 -1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_442
timestamp 1698431365
transform 1 0 5264 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_443
timestamp 1698431365
transform 1 0 13104 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_444
timestamp 1698431365
transform 1 0 20944 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_445
timestamp 1698431365
transform 1 0 28784 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_446
timestamp 1698431365
transform 1 0 36624 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_447
timestamp 1698431365
transform 1 0 44464 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_48_448
timestamp 1698431365
transform 1 0 52304 0 1 40768
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_449
timestamp 1698431365
transform 1 0 9184 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_450
timestamp 1698431365
transform 1 0 17024 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_451
timestamp 1698431365
transform 1 0 24864 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_452
timestamp 1698431365
transform 1 0 32704 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_453
timestamp 1698431365
transform 1 0 40544 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_49_454
timestamp 1698431365
transform 1 0 48384 0 -1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_455
timestamp 1698431365
transform 1 0 5264 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_456
timestamp 1698431365
transform 1 0 13104 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_457
timestamp 1698431365
transform 1 0 20944 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_458
timestamp 1698431365
transform 1 0 28784 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_459
timestamp 1698431365
transform 1 0 36624 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_460
timestamp 1698431365
transform 1 0 44464 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_50_461
timestamp 1698431365
transform 1 0 52304 0 1 42336
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_462
timestamp 1698431365
transform 1 0 9184 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_463
timestamp 1698431365
transform 1 0 17024 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_464
timestamp 1698431365
transform 1 0 24864 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_465
timestamp 1698431365
transform 1 0 32704 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_466
timestamp 1698431365
transform 1 0 40544 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_51_467
timestamp 1698431365
transform 1 0 48384 0 -1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_468
timestamp 1698431365
transform 1 0 5264 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_469
timestamp 1698431365
transform 1 0 13104 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_470
timestamp 1698431365
transform 1 0 20944 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_471
timestamp 1698431365
transform 1 0 28784 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_472
timestamp 1698431365
transform 1 0 36624 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_473
timestamp 1698431365
transform 1 0 44464 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_52_474
timestamp 1698431365
transform 1 0 52304 0 1 43904
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_475
timestamp 1698431365
transform 1 0 9184 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_476
timestamp 1698431365
transform 1 0 17024 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_477
timestamp 1698431365
transform 1 0 24864 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_478
timestamp 1698431365
transform 1 0 32704 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_479
timestamp 1698431365
transform 1 0 40544 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_53_480
timestamp 1698431365
transform 1 0 48384 0 -1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_481
timestamp 1698431365
transform 1 0 5264 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_482
timestamp 1698431365
transform 1 0 13104 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_483
timestamp 1698431365
transform 1 0 20944 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_484
timestamp 1698431365
transform 1 0 28784 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_485
timestamp 1698431365
transform 1 0 36624 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_486
timestamp 1698431365
transform 1 0 44464 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_54_487
timestamp 1698431365
transform 1 0 52304 0 1 45472
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_488
timestamp 1698431365
transform 1 0 9184 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_489
timestamp 1698431365
transform 1 0 17024 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_490
timestamp 1698431365
transform 1 0 24864 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_491
timestamp 1698431365
transform 1 0 32704 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_492
timestamp 1698431365
transform 1 0 40544 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_55_493
timestamp 1698431365
transform 1 0 48384 0 -1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_494
timestamp 1698431365
transform 1 0 5264 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_495
timestamp 1698431365
transform 1 0 13104 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_496
timestamp 1698431365
transform 1 0 20944 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_497
timestamp 1698431365
transform 1 0 28784 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_498
timestamp 1698431365
transform 1 0 36624 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_499
timestamp 1698431365
transform 1 0 44464 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_56_500
timestamp 1698431365
transform 1 0 52304 0 1 47040
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_501
timestamp 1698431365
transform 1 0 9184 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_502
timestamp 1698431365
transform 1 0 17024 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_503
timestamp 1698431365
transform 1 0 24864 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_504
timestamp 1698431365
transform 1 0 32704 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_505
timestamp 1698431365
transform 1 0 40544 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_57_506
timestamp 1698431365
transform 1 0 48384 0 -1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_507
timestamp 1698431365
transform 1 0 5264 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_508
timestamp 1698431365
transform 1 0 13104 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_509
timestamp 1698431365
transform 1 0 20944 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_510
timestamp 1698431365
transform 1 0 28784 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_511
timestamp 1698431365
transform 1 0 36624 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_512
timestamp 1698431365
transform 1 0 44464 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_58_513
timestamp 1698431365
transform 1 0 52304 0 1 48608
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_514
timestamp 1698431365
transform 1 0 9184 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_515
timestamp 1698431365
transform 1 0 17024 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_516
timestamp 1698431365
transform 1 0 24864 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_517
timestamp 1698431365
transform 1 0 32704 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_518
timestamp 1698431365
transform 1 0 40544 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_59_519
timestamp 1698431365
transform 1 0 48384 0 -1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_520
timestamp 1698431365
transform 1 0 5264 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_521
timestamp 1698431365
transform 1 0 13104 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_522
timestamp 1698431365
transform 1 0 20944 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_523
timestamp 1698431365
transform 1 0 28784 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_524
timestamp 1698431365
transform 1 0 36624 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_525
timestamp 1698431365
transform 1 0 44464 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_60_526
timestamp 1698431365
transform 1 0 52304 0 1 50176
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_527
timestamp 1698431365
transform 1 0 5152 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_528
timestamp 1698431365
transform 1 0 8960 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_529
timestamp 1698431365
transform 1 0 12768 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_530
timestamp 1698431365
transform 1 0 16576 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_531
timestamp 1698431365
transform 1 0 20384 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_532
timestamp 1698431365
transform 1 0 24192 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_533
timestamp 1698431365
transform 1 0 28000 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_534
timestamp 1698431365
transform 1 0 31808 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_535
timestamp 1698431365
transform 1 0 35616 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_536
timestamp 1698431365
transform 1 0 39424 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_537
timestamp 1698431365
transform 1 0 43232 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_538
timestamp 1698431365
transform 1 0 47040 0 -1 51744
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_61_539
timestamp 1698431365
transform 1 0 50848 0 -1 51744
box -86 -86 310 870
<< labels >>
flabel metal2 s 38528 0 38640 800 0 FreeSans 448 90 0 0 RXD
port 0 nsew signal input
flabel metal2 s 34048 0 34160 800 0 FreeSans 448 90 0 0 TXD
port 1 nsew signal tristate
flabel metal3 s 54200 3136 55000 3248 0 FreeSans 448 0 0 0 addr[0]
port 2 nsew signal input
flabel metal3 s 54200 5824 55000 5936 0 FreeSans 448 0 0 0 addr[1]
port 3 nsew signal input
flabel metal3 s 54200 8512 55000 8624 0 FreeSans 448 0 0 0 addr[2]
port 4 nsew signal input
flabel metal2 s 43008 0 43120 800 0 FreeSans 448 90 0 0 bus_cyc
port 5 nsew signal input
flabel metal2 s 47488 0 47600 800 0 FreeSans 448 90 0 0 bus_we
port 6 nsew signal input
flabel metal3 s 54200 11200 55000 11312 0 FreeSans 448 0 0 0 data_in[0]
port 7 nsew signal input
flabel metal3 s 54200 13888 55000 14000 0 FreeSans 448 0 0 0 data_in[1]
port 8 nsew signal input
flabel metal3 s 54200 16576 55000 16688 0 FreeSans 448 0 0 0 data_in[2]
port 9 nsew signal input
flabel metal3 s 54200 19264 55000 19376 0 FreeSans 448 0 0 0 data_in[3]
port 10 nsew signal input
flabel metal3 s 54200 21952 55000 22064 0 FreeSans 448 0 0 0 data_in[4]
port 11 nsew signal input
flabel metal3 s 54200 24640 55000 24752 0 FreeSans 448 0 0 0 data_in[5]
port 12 nsew signal input
flabel metal3 s 54200 27328 55000 27440 0 FreeSans 448 0 0 0 data_in[6]
port 13 nsew signal input
flabel metal3 s 54200 30016 55000 30128 0 FreeSans 448 0 0 0 data_in[7]
port 14 nsew signal input
flabel metal3 s 54200 32704 55000 32816 0 FreeSans 448 0 0 0 data_out[0]
port 15 nsew signal tristate
flabel metal3 s 54200 35392 55000 35504 0 FreeSans 448 0 0 0 data_out[1]
port 16 nsew signal tristate
flabel metal3 s 54200 38080 55000 38192 0 FreeSans 448 0 0 0 data_out[2]
port 17 nsew signal tristate
flabel metal3 s 54200 40768 55000 40880 0 FreeSans 448 0 0 0 data_out[3]
port 18 nsew signal tristate
flabel metal3 s 54200 43456 55000 43568 0 FreeSans 448 0 0 0 data_out[4]
port 19 nsew signal tristate
flabel metal3 s 54200 46144 55000 46256 0 FreeSans 448 0 0 0 data_out[5]
port 20 nsew signal tristate
flabel metal3 s 54200 48832 55000 48944 0 FreeSans 448 0 0 0 data_out[6]
port 21 nsew signal tristate
flabel metal3 s 54200 51520 55000 51632 0 FreeSans 448 0 0 0 data_out[7]
port 22 nsew signal tristate
flabel metal2 s 2688 0 2800 800 0 FreeSans 448 90 0 0 io_in
port 23 nsew signal input
flabel metal2 s 20608 0 20720 800 0 FreeSans 448 90 0 0 io_oeb[0]
port 24 nsew signal tristate
flabel metal2 s 25088 0 25200 800 0 FreeSans 448 90 0 0 io_oeb[1]
port 25 nsew signal tristate
flabel metal2 s 29568 0 29680 800 0 FreeSans 448 90 0 0 io_oeb[2]
port 26 nsew signal tristate
flabel metal2 s 7168 0 7280 800 0 FreeSans 448 90 0 0 io_out[0]
port 27 nsew signal tristate
flabel metal2 s 11648 0 11760 800 0 FreeSans 448 90 0 0 io_out[1]
port 28 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 io_out[2]
port 29 nsew signal tristate
flabel metal2 s 51968 0 52080 800 0 FreeSans 448 90 0 0 irq3
port 30 nsew signal tristate
flabel metal2 s 41216 54200 41328 55000 0 FreeSans 448 90 0 0 rst
port 31 nsew signal input
flabel metal4 s 4448 3076 4768 51804 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 35168 3076 35488 51804 0 FreeSans 1280 90 0 0 vdd
port 32 nsew power bidirectional
flabel metal4 s 19808 3076 20128 51804 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal4 s 50528 3076 50848 51804 0 FreeSans 1280 90 0 0 vss
port 33 nsew ground bidirectional
flabel metal2 s 13664 54200 13776 55000 0 FreeSans 448 90 0 0 wb_clk_i
port 34 nsew signal input
rlabel metal1 27496 50960 27496 50960 0 vdd
rlabel metal1 27496 51744 27496 51744 0 vss
rlabel metal2 38584 2086 38584 2086 0 RXD
rlabel metal2 34104 2198 34104 2198 0 TXD
rlabel metal2 45864 25928 45864 25928 0 _0000_
rlabel metal2 48832 28056 48832 28056 0 _0001_
rlabel metal2 51128 25872 51128 25872 0 _0002_
rlabel metal2 51128 22736 51128 22736 0 _0003_
rlabel metal2 51128 19656 51128 19656 0 _0004_
rlabel metal2 51128 17640 51128 17640 0 _0005_
rlabel metal2 50904 13384 50904 13384 0 _0006_
rlabel metal2 48888 12600 48888 12600 0 _0007_
rlabel metal2 50904 10248 50904 10248 0 _0008_
rlabel metal2 51128 7784 51128 7784 0 _0009_
rlabel metal3 50764 5768 50764 5768 0 _0010_
rlabel metal2 44968 4648 44968 4648 0 _0011_
rlabel metal2 41720 5264 41720 5264 0 _0012_
rlabel metal3 33544 4424 33544 4424 0 _0013_
rlabel metal2 42392 11760 42392 11760 0 _0014_
rlabel metal2 44520 15736 44520 15736 0 _0015_
rlabel metal2 41944 17696 41944 17696 0 _0016_
rlabel metal2 38136 11816 38136 11816 0 _0017_
rlabel metal3 35840 12040 35840 12040 0 _0018_
rlabel metal2 27944 14056 27944 14056 0 _0019_
rlabel metal3 30912 11480 30912 11480 0 _0020_
rlabel metal2 32424 8372 32424 8372 0 _0021_
rlabel metal2 39592 7784 39592 7784 0 _0022_
rlabel metal2 32536 6496 32536 6496 0 _0023_
rlabel metal2 27720 9352 27720 9352 0 _0024_
rlabel metal2 27048 12600 27048 12600 0 _0025_
rlabel metal2 22232 13328 22232 13328 0 _0026_
rlabel metal2 22176 11480 22176 11480 0 _0027_
rlabel metal2 21448 18032 21448 18032 0 _0028_
rlabel metal2 23464 15540 23464 15540 0 _0029_
rlabel metal2 24024 19600 24024 19600 0 _0030_
rlabel metal2 37688 4648 37688 4648 0 _0031_
rlabel metal3 35224 32424 35224 32424 0 _0032_
rlabel metal2 33208 33936 33208 33936 0 _0033_
rlabel metal2 30184 34160 30184 34160 0 _0034_
rlabel metal2 31080 34888 31080 34888 0 _0035_
rlabel metal2 30856 30464 30856 30464 0 _0036_
rlabel metal3 28896 28840 28896 28840 0 _0037_
rlabel metal3 28784 26152 28784 26152 0 _0038_
rlabel metal3 31248 27160 31248 27160 0 _0039_
rlabel metal3 49560 4424 49560 4424 0 _0040_
rlabel metal2 51128 29848 51128 29848 0 _0041_
rlabel metal2 45528 33712 45528 33712 0 _0042_
rlabel metal2 46312 36120 46312 36120 0 _0043_
rlabel metal2 51128 31304 51128 31304 0 _0044_
rlabel metal3 50512 33992 50512 33992 0 _0045_
rlabel metal2 51240 36848 51240 36848 0 _0046_
rlabel metal3 50512 41832 50512 41832 0 _0047_
rlabel metal2 51128 38976 51128 38976 0 _0048_
rlabel metal2 46536 50456 46536 50456 0 _0049_
rlabel metal2 51128 47152 51128 47152 0 _0050_
rlabel metal2 51240 49896 51240 49896 0 _0051_
rlabel metal2 50904 43876 50904 43876 0 _0052_
rlabel metal3 42000 29624 42000 29624 0 _0053_
rlabel metal2 26096 30856 26096 30856 0 _0054_
rlabel metal2 25816 34552 25816 34552 0 _0055_
rlabel metal2 22904 36120 22904 36120 0 _0056_
rlabel metal2 21448 33712 21448 33712 0 _0057_
rlabel metal2 20440 29736 20440 29736 0 _0058_
rlabel metal2 19712 26376 19712 26376 0 _0059_
rlabel metal2 19880 24024 19880 24024 0 _0060_
rlabel metal2 22512 23352 22512 23352 0 _0061_
rlabel metal2 36008 22064 36008 22064 0 _0062_
rlabel metal2 34328 24360 34328 24360 0 _0063_
rlabel metal3 35560 18424 35560 18424 0 _0064_
rlabel metal2 30744 18368 30744 18368 0 _0065_
rlabel metal3 28168 20440 28168 20440 0 _0066_
rlabel metal2 27944 22120 27944 22120 0 _0067_
rlabel metal2 31752 21168 31752 21168 0 _0068_
rlabel metal2 27048 18816 27048 18816 0 _0069_
rlabel metal2 29848 42280 29848 42280 0 _0070_
rlabel metal3 22624 40488 22624 40488 0 _0071_
rlabel metal2 26488 40712 26488 40712 0 _0072_
rlabel metal2 22344 39760 22344 39760 0 _0073_
rlabel metal3 22456 50456 22456 50456 0 _0074_
rlabel metal2 32648 50456 32648 50456 0 _0075_
rlabel metal3 29064 47320 29064 47320 0 _0076_
rlabel metal3 28000 50456 28000 50456 0 _0077_
rlabel metal2 33208 47768 33208 47768 0 _0078_
rlabel metal3 17080 50456 17080 50456 0 _0079_
rlabel metal2 16632 45136 16632 45136 0 _0080_
rlabel metal2 17080 42336 17080 42336 0 _0081_
rlabel metal3 10528 45304 10528 45304 0 _0082_
rlabel metal2 14280 48048 14280 48048 0 _0083_
rlabel metal2 9688 43120 9688 43120 0 _0084_
rlabel metal2 14280 40320 14280 40320 0 _0085_
rlabel metal2 38360 50456 38360 50456 0 _0086_
rlabel metal2 35112 49448 35112 49448 0 _0087_
rlabel metal2 42784 50456 42784 50456 0 _0088_
rlabel metal2 43064 47880 43064 47880 0 _0089_
rlabel metal2 44184 46312 44184 46312 0 _0090_
rlabel metal3 43904 44968 43904 44968 0 _0091_
rlabel metal2 41160 42392 41160 42392 0 _0092_
rlabel metal2 37128 46256 37128 46256 0 _0093_
rlabel metal2 29400 43960 29400 43960 0 _0094_
rlabel metal2 2296 15736 2296 15736 0 _0095_
rlabel metal2 2520 13328 2520 13328 0 _0096_
rlabel metal3 6664 18648 6664 18648 0 _0097_
rlabel metal2 2520 10920 2520 10920 0 _0098_
rlabel metal2 4760 9576 4760 9576 0 _0099_
rlabel metal2 7784 10360 7784 10360 0 _0100_
rlabel metal2 10696 9912 10696 9912 0 _0101_
rlabel metal2 12152 6776 12152 6776 0 _0102_
rlabel metal2 14392 10136 14392 10136 0 _0103_
rlabel metal2 17752 12096 17752 12096 0 _0104_
rlabel metal2 19320 17024 19320 17024 0 _0105_
rlabel metal2 16576 19096 16576 19096 0 _0106_
rlabel metal2 12600 17696 12600 17696 0 _0107_
rlabel metal2 10304 16744 10304 16744 0 _0108_
rlabel metal2 2520 23408 2520 23408 0 _0109_
rlabel metal2 2520 21896 2520 21896 0 _0110_
rlabel metal3 11256 23016 11256 23016 0 _0111_
rlabel metal2 11032 20552 11032 20552 0 _0112_
rlabel metal2 2520 26712 2520 26712 0 _0113_
rlabel metal2 2520 29064 2520 29064 0 _0114_
rlabel metal3 3976 32424 3976 32424 0 _0115_
rlabel metal3 4144 34776 4144 34776 0 _0116_
rlabel metal3 3808 37128 3808 37128 0 _0117_
rlabel metal2 5768 41216 5768 41216 0 _0118_
rlabel metal3 10080 39480 10080 39480 0 _0119_
rlabel metal3 11032 37240 11032 37240 0 _0120_
rlabel metal2 11480 29848 11480 29848 0 _0121_
rlabel metal2 10976 33096 10976 33096 0 _0122_
rlabel metal2 12712 28000 12712 28000 0 _0123_
rlabel metal2 11928 24864 11928 24864 0 _0124_
rlabel metal2 45640 32144 45640 32144 0 _0125_
rlabel metal2 9072 7672 9072 7672 0 _0126_
rlabel metal2 30072 4480 30072 4480 0 _0127_
rlabel metal2 26040 4648 26040 4648 0 _0128_
rlabel metal2 22400 4424 22400 4424 0 _0129_
rlabel metal2 18200 4816 18200 4816 0 _0130_
rlabel metal2 15288 5432 15288 5432 0 _0131_
rlabel metal2 16184 6720 16184 6720 0 _0132_
rlabel metal3 18816 8344 18816 8344 0 _0133_
rlabel metal2 23688 7728 23688 7728 0 _0134_
rlabel metal2 8568 7112 8568 7112 0 _0135_
rlabel metal2 38248 36848 38248 36848 0 _0136_
rlabel metal3 35728 41048 35728 41048 0 _0137_
rlabel metal3 35728 37912 35728 37912 0 _0138_
rlabel metal3 46592 40936 46592 40936 0 _0139_
rlabel metal2 44968 39144 44968 39144 0 _0140_
rlabel metal2 46984 39088 46984 39088 0 _0141_
rlabel metal3 44016 35784 44016 35784 0 _0142_
rlabel metal2 40600 39760 40600 39760 0 _0143_
rlabel metal2 10248 21056 10248 21056 0 _0144_
rlabel metal2 8120 25816 8120 25816 0 _0145_
rlabel metal2 7784 26040 7784 26040 0 _0146_
rlabel metal2 10416 21000 10416 21000 0 _0147_
rlabel metal3 7448 37240 7448 37240 0 _0148_
rlabel metal3 7168 29512 7168 29512 0 _0149_
rlabel metal2 6328 30352 6328 30352 0 _0150_
rlabel metal2 8344 22624 8344 22624 0 _0151_
rlabel metal2 5656 30128 5656 30128 0 _0152_
rlabel metal2 5544 27272 5544 27272 0 _0153_
rlabel metal2 9240 34944 9240 34944 0 _0154_
rlabel metal2 5544 26600 5544 26600 0 _0155_
rlabel metal2 6216 32200 6216 32200 0 _0156_
rlabel metal2 5208 29120 5208 29120 0 _0157_
rlabel metal2 2856 29064 2856 29064 0 _0158_
rlabel metal3 7728 31640 7728 31640 0 _0159_
rlabel metal2 5600 33208 5600 33208 0 _0160_
rlabel metal2 8232 28168 8232 28168 0 _0161_
rlabel metal2 5992 35000 5992 35000 0 _0162_
rlabel metal2 5712 32648 5712 32648 0 _0163_
rlabel metal2 6664 32760 6664 32760 0 _0164_
rlabel metal3 5712 32648 5712 32648 0 _0165_
rlabel metal2 5880 35168 5880 35168 0 _0166_
rlabel metal2 4984 34496 4984 34496 0 _0167_
rlabel metal2 5320 34440 5320 34440 0 _0168_
rlabel metal3 7224 38584 7224 38584 0 _0169_
rlabel metal2 7672 29400 7672 29400 0 _0170_
rlabel metal2 9016 34552 9016 34552 0 _0171_
rlabel metal2 7560 38724 7560 38724 0 _0172_
rlabel metal2 7224 39200 7224 39200 0 _0173_
rlabel metal2 5992 36624 5992 36624 0 _0174_
rlabel metal2 5320 37520 5320 37520 0 _0175_
rlabel metal2 6048 37464 6048 37464 0 _0176_
rlabel metal2 4872 37520 4872 37520 0 _0177_
rlabel metal3 5768 39480 5768 39480 0 _0178_
rlabel metal2 6552 40208 6552 40208 0 _0179_
rlabel metal2 5600 39480 5600 39480 0 _0180_
rlabel metal2 5992 40096 5992 40096 0 _0181_
rlabel metal2 8736 38248 8736 38248 0 _0182_
rlabel metal2 9576 37520 9576 37520 0 _0183_
rlabel metal2 10192 39032 10192 39032 0 _0184_
rlabel metal2 8568 38808 8568 38808 0 _0185_
rlabel metal2 9576 39704 9576 39704 0 _0186_
rlabel metal2 9464 37296 9464 37296 0 _0187_
rlabel metal2 10472 37576 10472 37576 0 _0188_
rlabel metal2 9912 37296 9912 37296 0 _0189_
rlabel metal3 40208 32648 40208 32648 0 _0190_
rlabel metal3 11648 30296 11648 30296 0 _0191_
rlabel metal2 9744 30968 9744 30968 0 _0192_
rlabel metal2 8960 35448 8960 35448 0 _0193_
rlabel metal2 10024 33320 10024 33320 0 _0194_
rlabel metal2 9352 31920 9352 31920 0 _0195_
rlabel metal2 9240 31304 9240 31304 0 _0196_
rlabel metal2 9912 30688 9912 30688 0 _0197_
rlabel metal2 11144 29232 11144 29232 0 _0198_
rlabel metal2 10920 33376 10920 33376 0 _0199_
rlabel metal2 9576 33040 9576 33040 0 _0200_
rlabel metal2 9912 32984 9912 32984 0 _0201_
rlabel metal2 9352 27832 9352 27832 0 _0202_
rlabel metal2 10304 28840 10304 28840 0 _0203_
rlabel metal2 10472 28000 10472 28000 0 _0204_
rlabel metal2 10248 27720 10248 27720 0 _0205_
rlabel metal2 10696 27384 10696 27384 0 _0206_
rlabel metal2 10808 25032 10808 25032 0 _0207_
rlabel metal2 9688 26152 9688 26152 0 _0208_
rlabel metal4 40040 40488 40040 40488 0 _0209_
rlabel metal2 38696 38668 38696 38668 0 _0210_
rlabel metal2 38920 31416 38920 31416 0 _0211_
rlabel metal2 39256 32144 39256 32144 0 _0212_
rlabel metal2 29176 4592 29176 4592 0 _0213_
rlabel metal2 29456 6664 29456 6664 0 _0214_
rlabel metal2 28168 5432 28168 5432 0 _0215_
rlabel metal2 18984 5488 18984 5488 0 _0216_
rlabel metal3 27216 5096 27216 5096 0 _0217_
rlabel metal2 20216 6664 20216 6664 0 _0218_
rlabel metal2 22680 5320 22680 5320 0 _0219_
rlabel metal3 20384 5320 20384 5320 0 _0220_
rlabel metal2 29064 7840 29064 7840 0 _0221_
rlabel metal2 19544 5656 19544 5656 0 _0222_
rlabel metal3 20328 7336 20328 7336 0 _0223_
rlabel metal3 20104 8120 20104 8120 0 _0224_
rlabel metal2 23352 7616 23352 7616 0 _0225_
rlabel metal2 8680 8176 8680 8176 0 _0226_
rlabel metal2 8120 7560 8120 7560 0 _0227_
rlabel metal2 39144 39984 39144 39984 0 _0228_
rlabel metal2 38696 37128 38696 37128 0 _0229_
rlabel metal2 37352 41832 37352 41832 0 _0230_
rlabel metal2 37072 39816 37072 39816 0 _0231_
rlabel metal2 45416 39424 45416 39424 0 _0232_
rlabel metal2 37408 38024 37408 38024 0 _0233_
rlabel metal2 36568 39004 36568 39004 0 _0234_
rlabel metal2 45416 42784 45416 42784 0 _0235_
rlabel metal2 45696 41160 45696 41160 0 _0236_
rlabel metal2 43960 40320 43960 40320 0 _0237_
rlabel metal2 44296 40824 44296 40824 0 _0238_
rlabel metal2 45192 41048 45192 41048 0 _0239_
rlabel metal2 44744 39480 44744 39480 0 _0240_
rlabel metal2 47096 39256 47096 39256 0 _0241_
rlabel metal2 46648 39088 46648 39088 0 _0242_
rlabel metal2 43288 39536 43288 39536 0 _0243_
rlabel metal2 43792 37352 43792 37352 0 _0244_
rlabel metal2 41160 40712 41160 40712 0 _0245_
rlabel metal2 40208 40152 40208 40152 0 _0246_
rlabel metal2 31192 9520 31192 9520 0 _0247_
rlabel metal2 18088 43792 18088 43792 0 _0248_
rlabel metal2 48888 9744 48888 9744 0 _0249_
rlabel metal2 38024 15344 38024 15344 0 _0250_
rlabel metal2 36568 16184 36568 16184 0 _0251_
rlabel metal2 33544 20860 33544 20860 0 _0252_
rlabel metal2 33544 17136 33544 17136 0 _0253_
rlabel metal2 34552 16184 34552 16184 0 _0254_
rlabel metal2 41048 10304 41048 10304 0 _0255_
rlabel metal2 45584 9800 45584 9800 0 _0256_
rlabel metal2 38584 16128 38584 16128 0 _0257_
rlabel metal3 37128 17416 37128 17416 0 _0258_
rlabel metal2 38136 16520 38136 16520 0 _0259_
rlabel metal2 32984 16688 32984 16688 0 _0260_
rlabel metal2 36344 16576 36344 16576 0 _0261_
rlabel metal2 38752 14504 38752 14504 0 _0262_
rlabel metal2 42056 17192 42056 17192 0 _0263_
rlabel metal3 39312 17640 39312 17640 0 _0264_
rlabel metal2 40040 16744 40040 16744 0 _0265_
rlabel metal2 38920 19096 38920 19096 0 _0266_
rlabel metal2 31192 19376 31192 19376 0 _0267_
rlabel metal2 38584 18368 38584 18368 0 _0268_
rlabel metal2 40488 15652 40488 15652 0 _0269_
rlabel metal2 41496 8624 41496 8624 0 _0270_
rlabel metal2 48552 10192 48552 10192 0 _0271_
rlabel metal3 46928 25480 46928 25480 0 _0272_
rlabel metal2 44800 20552 44800 20552 0 _0273_
rlabel metal2 43512 23016 43512 23016 0 _0274_
rlabel metal2 42840 23072 42840 23072 0 _0275_
rlabel metal2 43064 20384 43064 20384 0 _0276_
rlabel metal2 43624 22624 43624 22624 0 _0277_
rlabel metal2 31528 9688 31528 9688 0 _0278_
rlabel metal2 46648 11144 46648 11144 0 _0279_
rlabel metal2 26936 22064 26936 22064 0 _0280_
rlabel metal2 45752 24416 45752 24416 0 _0281_
rlabel metal2 46312 25200 46312 25200 0 _0282_
rlabel metal3 22904 22120 22904 22120 0 _0283_
rlabel metal2 41552 34888 41552 34888 0 _0284_
rlabel metal2 41496 40712 41496 40712 0 _0285_
rlabel metal2 43064 24304 43064 24304 0 _0286_
rlabel metal2 42392 19544 42392 19544 0 _0287_
rlabel metal2 50624 22232 50624 22232 0 _0288_
rlabel metal2 49280 24920 49280 24920 0 _0289_
rlabel metal2 48888 22344 48888 22344 0 _0290_
rlabel metal2 48944 22568 48944 22568 0 _0291_
rlabel metal2 50288 25368 50288 25368 0 _0292_
rlabel metal3 48664 25256 48664 25256 0 _0293_
rlabel metal2 48104 26068 48104 26068 0 _0294_
rlabel metal3 31920 21168 31920 21168 0 _0295_
rlabel metal2 45976 19600 45976 19600 0 _0296_
rlabel metal2 51240 23800 51240 23800 0 _0297_
rlabel metal2 49896 25200 49896 25200 0 _0298_
rlabel metal2 49112 23744 49112 23744 0 _0299_
rlabel metal2 49784 25648 49784 25648 0 _0300_
rlabel metal2 51016 25928 51016 25928 0 _0301_
rlabel metal3 50008 22232 50008 22232 0 _0302_
rlabel metal2 49112 22064 49112 22064 0 _0303_
rlabel metal2 49560 22512 49560 22512 0 _0304_
rlabel metal2 50904 22792 50904 22792 0 _0305_
rlabel metal2 50680 15232 50680 15232 0 _0306_
rlabel metal2 49224 18760 49224 18760 0 _0307_
rlabel metal2 49560 19600 49560 19600 0 _0308_
rlabel metal2 49784 20832 49784 20832 0 _0309_
rlabel metal2 48888 19544 48888 19544 0 _0310_
rlabel metal2 49728 19208 49728 19208 0 _0311_
rlabel metal3 50512 19096 50512 19096 0 _0312_
rlabel metal2 50120 17136 50120 17136 0 _0313_
rlabel metal2 46424 14784 46424 14784 0 _0314_
rlabel metal3 48944 17640 48944 17640 0 _0315_
rlabel metal2 49448 18088 49448 18088 0 _0316_
rlabel metal3 50624 18312 50624 18312 0 _0317_
rlabel metal2 38248 11536 38248 11536 0 _0318_
rlabel metal2 49896 15736 49896 15736 0 _0319_
rlabel metal2 50232 16240 50232 16240 0 _0320_
rlabel metal2 50120 15624 50120 15624 0 _0321_
rlabel metal2 50512 13160 50512 13160 0 _0322_
rlabel metal2 48664 15736 48664 15736 0 _0323_
rlabel metal2 48160 16072 48160 16072 0 _0324_
rlabel metal2 48552 15176 48552 15176 0 _0325_
rlabel metal2 48776 12656 48776 12656 0 _0326_
rlabel metal3 51548 6552 51548 6552 0 _0327_
rlabel metal2 43064 8736 43064 8736 0 _0328_
rlabel metal2 25816 9856 25816 9856 0 _0329_
rlabel metal3 46088 10584 46088 10584 0 _0330_
rlabel metal3 48216 10584 48216 10584 0 _0331_
rlabel metal2 36904 7168 36904 7168 0 _0332_
rlabel metal2 49336 10192 49336 10192 0 _0333_
rlabel metal3 51548 8008 51548 8008 0 _0334_
rlabel metal2 47992 9744 47992 9744 0 _0335_
rlabel metal2 48832 8232 48832 8232 0 _0336_
rlabel metal2 48720 8120 48720 8120 0 _0337_
rlabel metal3 49672 8064 49672 8064 0 _0338_
rlabel metal2 49112 6720 49112 6720 0 _0339_
rlabel metal2 42504 6272 42504 6272 0 _0340_
rlabel metal2 48104 7896 48104 7896 0 _0341_
rlabel metal3 49056 6664 49056 6664 0 _0342_
rlabel metal2 49896 6216 49896 6216 0 _0343_
rlabel metal3 41944 6552 41944 6552 0 _0344_
rlabel metal2 45808 7448 45808 7448 0 _0345_
rlabel metal2 44800 5208 44800 5208 0 _0346_
rlabel metal3 40824 29512 40824 29512 0 _0347_
rlabel metal3 41608 29960 41608 29960 0 _0348_
rlabel metal3 46144 21000 46144 21000 0 _0349_
rlabel metal2 39928 9352 39928 9352 0 _0350_
rlabel metal3 31920 14112 31920 14112 0 _0351_
rlabel metal2 42224 6888 42224 6888 0 _0352_
rlabel metal2 42840 6888 42840 6888 0 _0353_
rlabel metal2 42672 6104 42672 6104 0 _0354_
rlabel metal2 42840 8232 42840 8232 0 _0355_
rlabel metal2 25592 22008 25592 22008 0 _0356_
rlabel metal2 33320 6496 33320 6496 0 _0357_
rlabel metal3 28952 7560 28952 7560 0 _0358_
rlabel metal2 31752 6328 31752 6328 0 _0359_
rlabel metal3 34888 5880 34888 5880 0 _0360_
rlabel metal2 43512 15568 43512 15568 0 _0361_
rlabel metal2 36232 10192 36232 10192 0 _0362_
rlabel metal2 39704 14112 39704 14112 0 _0363_
rlabel metal2 32424 14224 32424 14224 0 _0364_
rlabel metal2 42056 12152 42056 12152 0 _0365_
rlabel metal2 32312 7168 32312 7168 0 _0366_
rlabel metal3 41888 15288 41888 15288 0 _0367_
rlabel metal3 44240 14280 44240 14280 0 _0368_
rlabel metal2 35672 13048 35672 13048 0 _0369_
rlabel metal2 42616 16240 42616 16240 0 _0370_
rlabel metal3 43512 15400 43512 15400 0 _0371_
rlabel metal3 32424 15624 32424 15624 0 _0372_
rlabel metal3 44072 15176 44072 15176 0 _0373_
rlabel metal2 40712 14784 40712 14784 0 _0374_
rlabel metal2 41832 15876 41832 15876 0 _0375_
rlabel metal3 37352 12712 37352 12712 0 _0376_
rlabel metal2 38920 12936 38920 12936 0 _0377_
rlabel metal2 38472 12152 38472 12152 0 _0378_
rlabel metal2 35672 15288 35672 15288 0 _0379_
rlabel metal2 36232 13272 36232 13272 0 _0380_
rlabel metal2 36344 12320 36344 12320 0 _0381_
rlabel metal2 31640 15176 31640 15176 0 _0382_
rlabel metal2 31864 14560 31864 14560 0 _0383_
rlabel metal3 33376 14728 33376 14728 0 _0384_
rlabel metal3 31808 14392 31808 14392 0 _0385_
rlabel metal2 31640 14728 31640 14728 0 _0386_
rlabel metal2 31752 11564 31752 11564 0 _0387_
rlabel metal2 35504 10024 35504 10024 0 _0388_
rlabel metal3 33208 9800 33208 9800 0 _0389_
rlabel metal2 32088 11256 32088 11256 0 _0390_
rlabel metal2 31528 11312 31528 11312 0 _0391_
rlabel metal3 33264 9688 33264 9688 0 _0392_
rlabel metal2 33432 9352 33432 9352 0 _0393_
rlabel metal2 30576 8232 30576 8232 0 _0394_
rlabel metal2 30072 7728 30072 7728 0 _0395_
rlabel metal2 29400 5432 29400 5432 0 _0396_
rlabel metal2 38248 7448 38248 7448 0 _0397_
rlabel metal2 38360 7952 38360 7952 0 _0398_
rlabel metal2 31696 5320 31696 5320 0 _0399_
rlabel metal3 34216 6776 34216 6776 0 _0400_
rlabel metal2 27832 8176 27832 8176 0 _0401_
rlabel metal2 25480 17752 25480 17752 0 _0402_
rlabel metal2 27608 12320 27608 12320 0 _0403_
rlabel metal2 27384 10080 27384 10080 0 _0404_
rlabel metal2 26824 9520 26824 9520 0 _0405_
rlabel metal2 27384 12040 27384 12040 0 _0406_
rlabel metal2 22792 9856 22792 9856 0 _0407_
rlabel metal2 21448 10864 21448 10864 0 _0408_
rlabel metal2 22456 12880 22456 12880 0 _0409_
rlabel metal2 21840 21784 21840 21784 0 _0410_
rlabel metal2 21896 19096 21896 19096 0 _0411_
rlabel metal2 20776 11480 20776 11480 0 _0412_
rlabel metal3 23128 12152 23128 12152 0 _0413_
rlabel metal2 22008 10892 22008 10892 0 _0414_
rlabel metal2 21448 17528 21448 17528 0 _0415_
rlabel metal2 23128 12096 23128 12096 0 _0416_
rlabel metal2 23296 16296 23296 16296 0 _0417_
rlabel metal2 25424 9240 25424 9240 0 _0418_
rlabel metal2 25144 18760 25144 18760 0 _0419_
rlabel metal3 25312 20104 25312 20104 0 _0420_
rlabel metal2 38808 5656 38808 5656 0 _0421_
rlabel metal2 37632 5096 37632 5096 0 _0422_
rlabel metal2 34888 21952 34888 21952 0 _0423_
rlabel metal2 26264 28672 26264 28672 0 _0424_
rlabel metal2 41384 23352 41384 23352 0 _0425_
rlabel metal2 41160 27608 41160 27608 0 _0426_
rlabel metal2 34776 31444 34776 31444 0 _0427_
rlabel metal3 30016 33320 30016 33320 0 _0428_
rlabel metal2 34664 32256 34664 32256 0 _0429_
rlabel metal2 35560 24136 35560 24136 0 _0430_
rlabel metal3 32200 29960 32200 29960 0 _0431_
rlabel metal2 32984 23744 32984 23744 0 _0432_
rlabel metal3 30856 26824 30856 26824 0 _0433_
rlabel metal2 31360 30072 31360 30072 0 _0434_
rlabel metal2 32816 32648 32816 32648 0 _0435_
rlabel metal2 33432 33208 33432 33208 0 _0436_
rlabel metal2 31472 23688 31472 23688 0 _0437_
rlabel metal2 30352 32312 30352 32312 0 _0438_
rlabel metal2 29736 33544 29736 33544 0 _0439_
rlabel metal3 31192 19152 31192 19152 0 _0440_
rlabel metal2 31136 32760 31136 32760 0 _0441_
rlabel metal2 30744 33712 30744 33712 0 _0442_
rlabel metal2 31024 26152 31024 26152 0 _0443_
rlabel metal2 30520 30128 30520 30128 0 _0444_
rlabel metal3 29456 26824 29456 26824 0 _0445_
rlabel metal2 30184 30072 30184 30072 0 _0446_
rlabel metal2 29848 26544 29848 26544 0 _0447_
rlabel metal2 30296 26600 30296 26600 0 _0448_
rlabel metal2 29848 27832 29848 27832 0 _0449_
rlabel metal2 30072 28616 30072 28616 0 _0450_
rlabel metal2 29736 25200 29736 25200 0 _0451_
rlabel metal2 29736 25984 29736 25984 0 _0452_
rlabel metal2 29456 26376 29456 26376 0 _0453_
rlabel metal2 31752 25648 31752 25648 0 _0454_
rlabel metal2 30856 25760 30856 25760 0 _0455_
rlabel metal2 30632 26684 30632 26684 0 _0456_
rlabel metal2 47656 10164 47656 10164 0 _0457_
rlabel metal2 42504 47432 42504 47432 0 _0458_
rlabel metal2 49784 33880 49784 33880 0 _0459_
rlabel metal2 47992 31248 47992 31248 0 _0460_
rlabel metal2 49056 37352 49056 37352 0 _0461_
rlabel metal2 36904 30632 36904 30632 0 _0462_
rlabel metal2 42336 25592 42336 25592 0 _0463_
rlabel via2 43400 33544 43400 33544 0 _0464_
rlabel metal3 39424 34104 39424 34104 0 _0465_
rlabel metal2 39200 31192 39200 31192 0 _0466_
rlabel metal2 37800 27832 37800 27832 0 _0467_
rlabel metal3 25592 26824 25592 26824 0 _0468_
rlabel metal2 37632 31528 37632 31528 0 _0469_
rlabel metal3 38528 30968 38528 30968 0 _0470_
rlabel metal3 44128 30744 44128 30744 0 _0471_
rlabel metal3 44464 31080 44464 31080 0 _0472_
rlabel metal3 42448 23016 42448 23016 0 _0473_
rlabel metal2 26936 23744 26936 23744 0 _0474_
rlabel metal2 28840 24640 28840 24640 0 _0475_
rlabel metal2 41720 22232 41720 22232 0 _0476_
rlabel metal2 40040 22008 40040 22008 0 _0477_
rlabel metal2 31416 24752 31416 24752 0 _0478_
rlabel metal2 37128 25536 37128 25536 0 _0479_
rlabel metal2 39424 23240 39424 23240 0 _0480_
rlabel metal2 45136 31080 45136 31080 0 _0481_
rlabel metal3 49784 30408 49784 30408 0 _0482_
rlabel metal2 39368 34888 39368 34888 0 _0483_
rlabel metal2 39480 33992 39480 33992 0 _0484_
rlabel metal2 38024 26208 38024 26208 0 _0485_
rlabel metal2 38976 26376 38976 26376 0 _0486_
rlabel metal3 38416 23800 38416 23800 0 _0487_
rlabel metal2 39200 23912 39200 23912 0 _0488_
rlabel metal3 43344 25144 43344 25144 0 _0489_
rlabel metal2 45976 33488 45976 33488 0 _0490_
rlabel metal3 42280 35672 42280 35672 0 _0491_
rlabel metal2 33544 25592 33544 25592 0 _0492_
rlabel metal3 39312 26040 39312 26040 0 _0493_
rlabel metal2 40040 26068 40040 26068 0 _0494_
rlabel metal2 50008 51296 50008 51296 0 _0495_
rlabel metal2 46816 35784 46816 35784 0 _0496_
rlabel metal2 50960 39368 50960 39368 0 _0497_
rlabel metal2 43568 31192 43568 31192 0 _0498_
rlabel metal2 23464 28168 23464 28168 0 _0499_
rlabel metal2 24360 31472 24360 31472 0 _0500_
rlabel metal3 43064 30912 43064 30912 0 _0501_
rlabel metal2 50008 31472 50008 31472 0 _0502_
rlabel metal2 50792 31752 50792 31752 0 _0503_
rlabel metal2 43456 32760 43456 32760 0 _0504_
rlabel metal3 24696 25368 24696 25368 0 _0505_
rlabel metal2 23912 30352 23912 30352 0 _0506_
rlabel metal3 35504 26600 35504 26600 0 _0507_
rlabel metal2 42952 32368 42952 32368 0 _0508_
rlabel metal2 49896 33040 49896 33040 0 _0509_
rlabel metal2 50232 33488 50232 33488 0 _0510_
rlabel metal2 43512 32032 43512 32032 0 _0511_
rlabel metal2 42392 31584 42392 31584 0 _0512_
rlabel metal2 43288 28560 43288 28560 0 _0513_
rlabel metal2 50120 35280 50120 35280 0 _0514_
rlabel metal3 50904 36344 50904 36344 0 _0515_
rlabel metal2 51016 46928 51016 46928 0 _0516_
rlabel metal2 42504 30184 42504 30184 0 _0517_
rlabel metal2 24696 27216 24696 27216 0 _0518_
rlabel metal3 36008 27160 36008 27160 0 _0519_
rlabel metal2 48384 40936 48384 40936 0 _0520_
rlabel metal2 49112 41496 49112 41496 0 _0521_
rlabel metal2 39816 30884 39816 30884 0 _0522_
rlabel metal3 31920 25648 31920 25648 0 _0523_
rlabel metal2 39928 27384 39928 27384 0 _0524_
rlabel metal3 49896 39368 49896 39368 0 _0525_
rlabel metal2 51128 39592 51128 39592 0 _0526_
rlabel metal2 33096 42336 33096 42336 0 _0527_
rlabel metal2 15960 37688 15960 37688 0 _0528_
rlabel metal3 18536 36568 18536 36568 0 _0529_
rlabel metal2 18424 37296 18424 37296 0 _0530_
rlabel metal2 18592 37352 18592 37352 0 _0531_
rlabel metal3 18984 38920 18984 38920 0 _0532_
rlabel metal3 19208 37912 19208 37912 0 _0533_
rlabel metal2 20216 38360 20216 38360 0 _0534_
rlabel metal2 19432 39060 19432 39060 0 _0535_
rlabel metal3 17976 38360 17976 38360 0 _0536_
rlabel metal2 19880 38724 19880 38724 0 _0537_
rlabel metal2 19544 40320 19544 40320 0 _0538_
rlabel metal2 32424 39592 32424 39592 0 _0539_
rlabel metal2 32928 38808 32928 38808 0 _0540_
rlabel metal2 30688 38808 30688 38808 0 _0541_
rlabel metal2 30968 38780 30968 38780 0 _0542_
rlabel metal2 32088 38304 32088 38304 0 _0543_
rlabel metal2 29512 37632 29512 37632 0 _0544_
rlabel metal3 27608 37240 27608 37240 0 _0545_
rlabel metal2 28560 36568 28560 36568 0 _0546_
rlabel metal2 26488 37744 26488 37744 0 _0547_
rlabel metal2 31976 37688 31976 37688 0 _0548_
rlabel metal2 33208 41664 33208 41664 0 _0549_
rlabel metal2 47544 44240 47544 44240 0 _0550_
rlabel metal2 49336 48160 49336 48160 0 _0551_
rlabel metal2 34888 44688 34888 44688 0 _0552_
rlabel metal2 38808 45192 38808 45192 0 _0553_
rlabel metal3 44800 45192 44800 45192 0 _0554_
rlabel metal2 47096 48720 47096 48720 0 _0555_
rlabel metal2 49672 47376 49672 47376 0 _0556_
rlabel metal2 50624 47320 50624 47320 0 _0557_
rlabel metal2 50456 50680 50456 50680 0 _0558_
rlabel metal3 50176 51352 50176 51352 0 _0559_
rlabel metal2 51688 51632 51688 51632 0 _0560_
rlabel metal2 50008 45472 50008 45472 0 _0561_
rlabel metal2 49000 44464 49000 44464 0 _0562_
rlabel metal2 48272 45192 48272 45192 0 _0563_
rlabel metal2 48552 44520 48552 44520 0 _0564_
rlabel metal2 49392 43512 49392 43512 0 _0565_
rlabel metal2 49672 43904 49672 43904 0 _0566_
rlabel metal2 32200 24808 32200 24808 0 _0567_
rlabel metal2 38304 29512 38304 29512 0 _0568_
rlabel metal2 39368 29400 39368 29400 0 _0569_
rlabel metal2 23464 31808 23464 31808 0 _0570_
rlabel metal2 25592 33040 25592 33040 0 _0571_
rlabel metal2 25592 31696 25592 31696 0 _0572_
rlabel metal2 19096 20496 19096 20496 0 _0573_
rlabel metal2 12152 10752 12152 10752 0 _0574_
rlabel metal2 25928 33712 25928 33712 0 _0575_
rlabel metal3 19712 25480 19712 25480 0 _0576_
rlabel metal2 22232 35280 22232 35280 0 _0577_
rlabel metal2 25480 34384 25480 34384 0 _0578_
rlabel metal2 23184 33320 23184 33320 0 _0579_
rlabel metal2 22624 35784 22624 35784 0 _0580_
rlabel metal2 22792 32984 22792 32984 0 _0581_
rlabel metal2 21056 33320 21056 33320 0 _0582_
rlabel metal2 20104 24192 20104 24192 0 _0583_
rlabel metal2 20328 29064 20328 29064 0 _0584_
rlabel metal2 20664 28952 20664 28952 0 _0585_
rlabel metal2 21056 30184 21056 30184 0 _0586_
rlabel metal3 19544 27048 19544 27048 0 _0587_
rlabel metal2 19712 27048 19712 27048 0 _0588_
rlabel metal3 20104 24696 20104 24696 0 _0589_
rlabel metal2 19544 25032 19544 25032 0 _0590_
rlabel metal2 22680 23912 22680 23912 0 _0591_
rlabel metal2 22344 23800 22344 23800 0 _0592_
rlabel metal2 27720 21952 27720 21952 0 _0593_
rlabel metal2 31304 24192 31304 24192 0 _0594_
rlabel metal2 30632 21224 30632 21224 0 _0595_
rlabel metal2 29512 21504 29512 21504 0 _0596_
rlabel metal3 36400 22232 36400 22232 0 _0597_
rlabel metal2 31808 23912 31808 23912 0 _0598_
rlabel metal2 33208 24304 33208 24304 0 _0599_
rlabel metal2 34216 24192 34216 24192 0 _0600_
rlabel metal2 34552 23800 34552 23800 0 _0601_
rlabel metal3 34944 19096 34944 19096 0 _0602_
rlabel metal3 29792 23352 29792 23352 0 _0603_
rlabel metal3 32368 19096 32368 19096 0 _0604_
rlabel metal2 28336 20216 28336 20216 0 _0605_
rlabel metal3 29400 20776 29400 20776 0 _0606_
rlabel metal2 27944 22736 27944 22736 0 _0607_
rlabel metal3 28728 22344 28728 22344 0 _0608_
rlabel metal2 33992 21672 33992 21672 0 _0609_
rlabel metal3 27888 20104 27888 20104 0 _0610_
rlabel metal2 27720 20720 27720 20720 0 _0611_
rlabel metal2 26824 42056 26824 42056 0 _0612_
rlabel metal2 19768 44800 19768 44800 0 _0613_
rlabel metal2 26040 43680 26040 43680 0 _0614_
rlabel metal3 35224 45080 35224 45080 0 _0615_
rlabel metal2 34216 45416 34216 45416 0 _0616_
rlabel metal3 19992 44968 19992 44968 0 _0617_
rlabel metal3 23968 48328 23968 48328 0 _0618_
rlabel metal2 26824 43652 26824 43652 0 _0619_
rlabel metal2 29736 43176 29736 43176 0 _0620_
rlabel metal2 23800 42448 23800 42448 0 _0621_
rlabel metal2 25480 44408 25480 44408 0 _0622_
rlabel metal2 26264 43736 26264 43736 0 _0623_
rlabel metal2 33656 45248 33656 45248 0 _0624_
rlabel metal2 23464 44968 23464 44968 0 _0625_
rlabel metal2 25256 49392 25256 49392 0 _0626_
rlabel metal2 25816 43848 25816 43848 0 _0627_
rlabel metal2 20944 43624 20944 43624 0 _0628_
rlabel metal3 24584 50512 24584 50512 0 _0629_
rlabel metal2 26040 41216 26040 41216 0 _0630_
rlabel metal2 16352 44184 16352 44184 0 _0631_
rlabel metal2 23632 42168 23632 42168 0 _0632_
rlabel metal3 20496 44184 20496 44184 0 _0633_
rlabel metal3 25144 41160 25144 41160 0 _0634_
rlabel metal2 26544 41384 26544 41384 0 _0635_
rlabel metal2 23912 40600 23912 40600 0 _0636_
rlabel metal3 23968 40376 23968 40376 0 _0637_
rlabel metal2 22008 44072 22008 44072 0 _0638_
rlabel metal2 22680 45304 22680 45304 0 _0639_
rlabel metal2 22904 45360 22904 45360 0 _0640_
rlabel metal2 23072 40488 23072 40488 0 _0641_
rlabel metal2 20664 22512 20664 22512 0 _0642_
rlabel metal2 23464 46312 23464 46312 0 _0643_
rlabel metal2 26040 47488 26040 47488 0 _0644_
rlabel metal3 22904 48216 22904 48216 0 _0645_
rlabel metal3 25536 50456 25536 50456 0 _0646_
rlabel metal2 24360 50624 24360 50624 0 _0647_
rlabel metal2 20664 47712 20664 47712 0 _0648_
rlabel metal2 24080 50008 24080 50008 0 _0649_
rlabel metal2 39816 48776 39816 48776 0 _0650_
rlabel metal2 25704 49224 25704 49224 0 _0651_
rlabel metal2 24584 49056 24584 49056 0 _0652_
rlabel metal3 28672 49672 28672 49672 0 _0653_
rlabel metal2 26600 48720 26600 48720 0 _0654_
rlabel metal2 27048 48720 27048 48720 0 _0655_
rlabel metal2 27776 46872 27776 46872 0 _0656_
rlabel metal2 25704 47488 25704 47488 0 _0657_
rlabel metal3 27328 47432 27328 47432 0 _0658_
rlabel metal2 27608 50232 27608 50232 0 _0659_
rlabel metal2 26992 49224 26992 49224 0 _0660_
rlabel metal2 26992 50568 26992 50568 0 _0661_
rlabel metal2 22568 46592 22568 46592 0 _0662_
rlabel metal2 21336 47768 21336 47768 0 _0663_
rlabel metal2 19432 46984 19432 46984 0 _0664_
rlabel metal3 21280 48328 21280 48328 0 _0665_
rlabel metal2 21112 48160 21112 48160 0 _0666_
rlabel metal3 20048 48440 20048 48440 0 _0667_
rlabel metal3 26544 48104 26544 48104 0 _0668_
rlabel metal2 18424 49392 18424 49392 0 _0669_
rlabel metal2 18200 49168 18200 49168 0 _0670_
rlabel metal3 19824 48776 19824 48776 0 _0671_
rlabel metal2 19320 49504 19320 49504 0 _0672_
rlabel metal2 17416 48608 17416 48608 0 _0673_
rlabel metal2 18984 45304 18984 45304 0 _0674_
rlabel metal2 17640 44576 17640 44576 0 _0675_
rlabel metal2 19880 44576 19880 44576 0 _0676_
rlabel metal3 18200 44408 18200 44408 0 _0677_
rlabel metal3 19936 44072 19936 44072 0 _0678_
rlabel metal2 20104 43680 20104 43680 0 _0679_
rlabel metal3 19712 43512 19712 43512 0 _0680_
rlabel metal3 20720 46760 20720 46760 0 _0681_
rlabel metal3 18116 46872 18116 46872 0 _0682_
rlabel metal2 14504 46200 14504 46200 0 _0683_
rlabel metal2 13160 46312 13160 46312 0 _0684_
rlabel metal2 11648 45080 11648 45080 0 _0685_
rlabel metal3 11984 45192 11984 45192 0 _0686_
rlabel metal2 13272 47096 13272 47096 0 _0687_
rlabel metal2 14896 46648 14896 46648 0 _0688_
rlabel metal2 14672 47432 14672 47432 0 _0689_
rlabel metal2 12656 42168 12656 42168 0 _0690_
rlabel metal2 14056 43008 14056 43008 0 _0691_
rlabel metal2 14392 43232 14392 43232 0 _0692_
rlabel metal2 14728 43120 14728 43120 0 _0693_
rlabel metal3 12936 43624 12936 43624 0 _0694_
rlabel metal2 12376 43568 12376 43568 0 _0695_
rlabel metal2 15400 41664 15400 41664 0 _0696_
rlabel metal2 14392 41440 14392 41440 0 _0697_
rlabel metal3 15148 42504 15148 42504 0 _0698_
rlabel metal3 43736 42952 43736 42952 0 _0699_
rlabel metal2 36960 45752 36960 45752 0 _0700_
rlabel metal2 40264 46256 40264 46256 0 _0701_
rlabel metal2 40040 47936 40040 47936 0 _0702_
rlabel metal2 39816 45752 39816 45752 0 _0703_
rlabel metal2 38696 47880 38696 47880 0 _0704_
rlabel metal2 38360 49336 38360 49336 0 _0705_
rlabel metal2 35504 49224 35504 49224 0 _0706_
rlabel metal2 42112 48440 42112 48440 0 _0707_
rlabel metal2 41272 49336 41272 49336 0 _0708_
rlabel metal2 42056 46536 42056 46536 0 _0709_
rlabel metal3 42336 47320 42336 47320 0 _0710_
rlabel metal3 43512 45752 43512 45752 0 _0711_
rlabel metal2 42952 45248 42952 45248 0 _0712_
rlabel metal2 2632 28560 2632 28560 0 _0713_
rlabel metal2 41272 43456 41272 43456 0 _0714_
rlabel metal3 38724 46536 38724 46536 0 _0715_
rlabel metal3 35840 42168 35840 42168 0 _0716_
rlabel metal3 41608 42616 41608 42616 0 _0717_
rlabel metal2 38808 43120 38808 43120 0 _0718_
rlabel metal2 10696 24752 10696 24752 0 _0719_
rlabel metal2 16856 25088 16856 25088 0 _0720_
rlabel metal2 19096 24808 19096 24808 0 _0721_
rlabel metal2 15848 34216 15848 34216 0 _0722_
rlabel metal2 16296 30576 16296 30576 0 _0723_
rlabel metal2 16296 27720 16296 27720 0 _0724_
rlabel metal2 18424 28616 18424 28616 0 _0725_
rlabel metal3 18144 27720 18144 27720 0 _0726_
rlabel metal2 17416 28168 17416 28168 0 _0727_
rlabel metal2 15512 28616 15512 28616 0 _0728_
rlabel metal3 17752 28056 17752 28056 0 _0729_
rlabel metal2 17080 22512 17080 22512 0 _0730_
rlabel metal2 7112 20048 7112 20048 0 _0731_
rlabel metal2 20440 33096 20440 33096 0 _0732_
rlabel metal2 19544 32872 19544 32872 0 _0733_
rlabel metal2 18704 32536 18704 32536 0 _0734_
rlabel metal2 18816 31080 18816 31080 0 _0735_
rlabel metal3 17640 32648 17640 32648 0 _0736_
rlabel metal2 15512 32872 15512 32872 0 _0737_
rlabel metal2 15232 32536 15232 32536 0 _0738_
rlabel metal2 15008 32536 15008 32536 0 _0739_
rlabel metal3 14616 32536 14616 32536 0 _0740_
rlabel metal2 15848 32536 15848 32536 0 _0741_
rlabel metal3 16520 19992 16520 19992 0 _0742_
rlabel metal2 7616 19096 7616 19096 0 _0743_
rlabel metal3 7280 13160 7280 13160 0 _0744_
rlabel metal3 40712 21560 40712 21560 0 _0745_
rlabel metal2 10080 13944 10080 13944 0 _0746_
rlabel metal2 8568 15792 8568 15792 0 _0747_
rlabel metal2 8232 15456 8232 15456 0 _0748_
rlabel metal2 5096 18088 5096 18088 0 _0749_
rlabel metal2 5096 14364 5096 14364 0 _0750_
rlabel metal3 8344 18984 8344 18984 0 _0751_
rlabel metal3 12264 19096 12264 19096 0 _0752_
rlabel metal2 14168 20832 14168 20832 0 _0753_
rlabel metal2 7672 17304 7672 17304 0 _0754_
rlabel metal2 7392 15064 7392 15064 0 _0755_
rlabel metal3 5096 15288 5096 15288 0 _0756_
rlabel metal2 5992 13328 5992 13328 0 _0757_
rlabel metal2 16632 19824 16632 19824 0 _0758_
rlabel metal2 10472 14784 10472 14784 0 _0759_
rlabel metal2 7224 13888 7224 13888 0 _0760_
rlabel metal2 6776 14504 6776 14504 0 _0761_
rlabel metal2 6216 14000 6216 14000 0 _0762_
rlabel metal2 6888 13216 6888 13216 0 _0763_
rlabel metal2 7896 8316 7896 8316 0 _0764_
rlabel metal2 30520 5208 30520 5208 0 _0765_
rlabel metal2 6160 18424 6160 18424 0 _0766_
rlabel metal2 6664 18536 6664 18536 0 _0767_
rlabel metal2 5880 11872 5880 11872 0 _0768_
rlabel metal2 6552 18424 6552 18424 0 _0769_
rlabel metal2 5376 11256 5376 11256 0 _0770_
rlabel metal2 6328 12040 6328 12040 0 _0771_
rlabel metal2 12376 16184 12376 16184 0 _0772_
rlabel metal2 12096 14504 12096 14504 0 _0773_
rlabel metal2 10976 11256 10976 11256 0 _0774_
rlabel metal2 8568 11200 8568 11200 0 _0775_
rlabel metal2 7336 10640 7336 10640 0 _0776_
rlabel metal3 11480 11928 11480 11928 0 _0777_
rlabel metal2 8792 11648 8792 11648 0 _0778_
rlabel metal3 6944 11480 6944 11480 0 _0779_
rlabel metal2 13328 9240 13328 9240 0 _0780_
rlabel metal2 12824 10976 12824 10976 0 _0781_
rlabel metal2 10752 12152 10752 12152 0 _0782_
rlabel metal2 10976 10360 10976 10360 0 _0783_
rlabel metal3 13272 10584 13272 10584 0 _0784_
rlabel metal2 14840 12824 14840 12824 0 _0785_
rlabel metal2 12936 12096 12936 12096 0 _0786_
rlabel metal2 12264 11200 12264 11200 0 _0787_
rlabel metal2 14392 11480 14392 11480 0 _0788_
rlabel metal2 14392 14280 14392 14280 0 _0789_
rlabel metal2 14056 12432 14056 12432 0 _0790_
rlabel metal2 14616 11480 14616 11480 0 _0791_
rlabel metal3 17360 11368 17360 11368 0 _0792_
rlabel metal3 17248 11928 17248 11928 0 _0793_
rlabel metal2 18424 15204 18424 15204 0 _0794_
rlabel metal2 15848 13440 15848 13440 0 _0795_
rlabel metal2 15624 12768 15624 12768 0 _0796_
rlabel metal3 19880 14504 19880 14504 0 _0797_
rlabel metal3 17752 16856 17752 16856 0 _0798_
rlabel metal3 16520 15960 16520 15960 0 _0799_
rlabel metal3 19320 13608 19320 13608 0 _0800_
rlabel metal2 18648 13552 18648 13552 0 _0801_
rlabel metal2 17752 17528 17752 17528 0 _0802_
rlabel metal2 19096 15008 19096 15008 0 _0803_
rlabel metal3 18200 16632 18200 16632 0 _0804_
rlabel metal2 16072 17024 16072 17024 0 _0805_
rlabel metal3 16912 16072 16912 16072 0 _0806_
rlabel metal2 16408 16240 16408 16240 0 _0807_
rlabel metal2 16688 16856 16688 16856 0 _0808_
rlabel metal2 11704 16632 11704 16632 0 _0809_
rlabel metal2 15288 16576 15288 16576 0 _0810_
rlabel metal3 13944 16856 13944 16856 0 _0811_
rlabel metal2 5880 23632 5880 23632 0 _0812_
rlabel metal2 6440 19936 6440 19936 0 _0813_
rlabel metal2 10248 23072 10248 23072 0 _0814_
rlabel metal2 10584 23912 10584 23912 0 _0815_
rlabel metal2 6888 21952 6888 21952 0 _0816_
rlabel metal2 5768 23968 5768 23968 0 _0817_
rlabel metal2 2856 23464 2856 23464 0 _0818_
rlabel metal2 7672 23296 7672 23296 0 _0819_
rlabel metal2 5824 22344 5824 22344 0 _0820_
rlabel metal3 5600 23240 5600 23240 0 _0821_
rlabel metal3 6888 25256 6888 25256 0 _0822_
rlabel metal2 6104 24752 6104 24752 0 _0823_
rlabel metal2 5656 22624 5656 22624 0 _0824_
rlabel metal3 15260 23800 15260 23800 0 _0825_
rlabel metal2 9128 22456 9128 22456 0 _0826_
rlabel metal2 9352 23520 9352 23520 0 _0827_
rlabel metal2 8680 23576 8680 23576 0 _0828_
rlabel metal2 8456 23072 8456 23072 0 _0829_
rlabel metal2 53256 3304 53256 3304 0 addr[0]
rlabel metal2 52024 6272 52024 6272 0 addr[1]
rlabel metal2 53256 8792 53256 8792 0 addr[2]
rlabel metal2 43400 3416 43400 3416 0 bus_cyc
rlabel metal2 47544 2058 47544 2058 0 bus_we
rlabel metal2 37968 22456 37968 22456 0 clknet_0_wb_clk_i
rlabel metal2 1848 11760 1848 11760 0 clknet_4_0_0_wb_clk_i
rlabel metal2 50456 19320 50456 19320 0 clknet_4_10_0_wb_clk_i
rlabel metal2 50456 24696 50456 24696 0 clknet_4_11_0_wb_clk_i
rlabel metal3 33152 35336 33152 35336 0 clknet_4_12_0_wb_clk_i
rlabel metal2 34048 50568 34048 50568 0 clknet_4_13_0_wb_clk_i
rlabel metal2 49672 39200 49672 39200 0 clknet_4_14_0_wb_clk_i
rlabel metal2 45248 50456 45248 50456 0 clknet_4_15_0_wb_clk_i
rlabel metal2 1848 16464 1848 16464 0 clknet_4_1_0_wb_clk_i
rlabel metal2 29288 3976 29288 3976 0 clknet_4_2_0_wb_clk_i
rlabel metal2 30968 20468 30968 20468 0 clknet_4_3_0_wb_clk_i
rlabel metal2 1848 22568 1848 22568 0 clknet_4_4_0_wb_clk_i
rlabel metal2 1736 31892 1736 31892 0 clknet_4_5_0_wb_clk_i
rlabel metal2 19152 26264 19152 26264 0 clknet_4_6_0_wb_clk_i
rlabel metal2 16688 40376 16688 40376 0 clknet_4_7_0_wb_clk_i
rlabel metal2 32984 5488 32984 5488 0 clknet_4_8_0_wb_clk_i
rlabel metal2 28840 26432 28840 26432 0 clknet_4_9_0_wb_clk_i
rlabel metal3 53746 11256 53746 11256 0 data_in[0]
rlabel metal2 53256 14112 53256 14112 0 data_in[1]
rlabel metal2 53144 16352 53144 16352 0 data_in[2]
rlabel metal2 53256 19264 53256 19264 0 data_in[3]
rlabel metal2 53368 21896 53368 21896 0 data_in[4]
rlabel metal3 53746 24696 53746 24696 0 data_in[5]
rlabel metal2 53256 27608 53256 27608 0 data_in[6]
rlabel metal3 53746 30072 53746 30072 0 data_in[7]
rlabel metal2 53032 32592 53032 32592 0 data_out[0]
rlabel metal3 53634 35448 53634 35448 0 data_out[1]
rlabel metal3 53634 38136 53634 38136 0 data_out[2]
rlabel metal2 51912 41048 51912 41048 0 data_out[3]
rlabel metal3 53634 43512 53634 43512 0 data_out[4]
rlabel metal2 53032 47096 53032 47096 0 data_out[5]
rlabel metal2 51912 49000 51912 49000 0 data_out[6]
rlabel metal3 52682 51576 52682 51576 0 data_out[7]
rlabel metal2 2744 2086 2744 2086 0 io_in
rlabel metal2 7224 2086 7224 2086 0 io_out[0]
rlabel metal2 11704 2422 11704 2422 0 io_out[1]
rlabel metal2 52024 2198 52024 2198 0 irq3
rlabel metal3 39144 44072 39144 44072 0 net1
rlabel metal2 52920 19936 52920 19936 0 net10
rlabel metal2 52920 21952 52920 21952 0 net11
rlabel metal2 52920 24584 52920 24584 0 net12
rlabel metal3 48552 23688 48552 23688 0 net13
rlabel metal3 48328 17416 48328 17416 0 net14
rlabel metal2 3304 3808 3304 3808 0 net15
rlabel metal2 41216 50904 41216 50904 0 net16
rlabel metal2 10808 4984 10808 4984 0 net17
rlabel metal2 49448 31528 49448 31528 0 net18
rlabel metal2 49336 34496 49336 34496 0 net19
rlabel metal2 52696 4312 52696 4312 0 net2
rlabel metal2 50680 39872 50680 39872 0 net20
rlabel metal2 50008 39900 50008 39900 0 net21
rlabel metal2 51128 44744 51128 44744 0 net22
rlabel metal2 51184 48216 51184 48216 0 net23
rlabel metal2 53256 41496 53256 41496 0 net24
rlabel metal2 51128 44296 51128 44296 0 net25
rlabel metal2 11928 3584 11928 3584 0 net26
rlabel metal2 14392 4368 14392 4368 0 net27
rlabel metal2 48776 3864 48776 3864 0 net28
rlabel metal2 20664 2030 20664 2030 0 net29
rlabel metal2 51576 6384 51576 6384 0 net3
rlabel metal2 25144 2030 25144 2030 0 net30
rlabel metal2 16184 2030 16184 2030 0 net31
rlabel metal2 29624 2198 29624 2198 0 net32
rlabel metal2 52920 9632 52920 9632 0 net4
rlabel metal2 44968 21392 44968 21392 0 net5
rlabel metal2 45360 21448 45360 21448 0 net6
rlabel metal2 52920 11648 52920 11648 0 net7
rlabel metal3 12992 12152 12992 12152 0 net8
rlabel metal2 52864 15960 52864 15960 0 net9
rlabel metal2 41272 52906 41272 52906 0 rst
rlabel metal2 36232 5936 36232 5936 0 spi.busy
rlabel metal2 53312 6776 53312 6776 0 spi.counter\[0\]
rlabel metal2 53256 7672 53256 7672 0 spi.counter\[1\]
rlabel metal2 53256 5432 53256 5432 0 spi.counter\[2\]
rlabel metal3 46480 6552 46480 6552 0 spi.counter\[3\]
rlabel metal2 46312 5880 46312 5880 0 spi.counter\[4\]
rlabel metal2 31640 5040 31640 5040 0 spi.data_in_buff\[0\]
rlabel metal2 27608 6328 27608 6328 0 spi.data_in_buff\[1\]
rlabel metal2 22904 6216 22904 6216 0 spi.data_in_buff\[2\]
rlabel metal2 21336 7728 21336 7728 0 spi.data_in_buff\[3\]
rlabel metal2 20160 7672 20160 7672 0 spi.data_in_buff\[4\]
rlabel metal3 21280 8232 21280 8232 0 spi.data_in_buff\[5\]
rlabel via2 22232 8904 22232 8904 0 spi.data_in_buff\[6\]
rlabel metal2 25928 8288 25928 8288 0 spi.data_in_buff\[7\]
rlabel metal3 47208 25368 47208 25368 0 spi.data_out_buff\[0\]
rlabel metal2 49672 26096 49672 26096 0 spi.data_out_buff\[1\]
rlabel metal2 53256 25872 53256 25872 0 spi.data_out_buff\[2\]
rlabel metal2 50456 22344 50456 22344 0 spi.data_out_buff\[3\]
rlabel metal2 50120 19208 50120 19208 0 spi.data_out_buff\[4\]
rlabel metal3 50792 16688 50792 16688 0 spi.data_out_buff\[5\]
rlabel metal3 49280 14504 49280 14504 0 spi.data_out_buff\[6\]
rlabel metal2 46872 13160 46872 13160 0 spi.data_out_buff\[7\]
rlabel metal2 38024 16856 38024 16856 0 spi.div_counter\[0\]
rlabel metal2 38304 15960 38304 15960 0 spi.div_counter\[1\]
rlabel metal2 43288 17976 43288 17976 0 spi.div_counter\[2\]
rlabel metal2 34776 16688 34776 16688 0 spi.div_counter\[3\]
rlabel metal3 34496 12712 34496 12712 0 spi.div_counter\[4\]
rlabel metal2 30800 15288 30800 15288 0 spi.div_counter\[5\]
rlabel metal2 32872 16520 32872 16520 0 spi.div_counter\[6\]
rlabel metal2 34608 9688 34608 9688 0 spi.div_counter\[7\]
rlabel metal2 37128 21784 37128 21784 0 spi.divisor\[0\]
rlabel metal2 36680 24528 36680 24528 0 spi.divisor\[1\]
rlabel metal2 38360 18592 38360 18592 0 spi.divisor\[2\]
rlabel metal2 34888 26264 34888 26264 0 spi.divisor\[3\]
rlabel metal3 30296 20216 30296 20216 0 spi.divisor\[4\]
rlabel metal2 29400 22624 29400 22624 0 spi.divisor\[5\]
rlabel metal2 33824 20888 33824 20888 0 spi.divisor\[6\]
rlabel metal2 29904 20888 29904 20888 0 spi.divisor\[7\]
rlabel metal2 35784 6664 35784 6664 0 spi.dout\[0\]
rlabel metal2 27944 10864 27944 10864 0 spi.dout\[1\]
rlabel metal2 28784 24920 28784 24920 0 spi.dout\[2\]
rlabel metal2 24360 14364 24360 14364 0 spi.dout\[3\]
rlabel metal2 24136 12488 24136 12488 0 spi.dout\[4\]
rlabel metal2 22792 18704 22792 18704 0 spi.dout\[5\]
rlabel metal2 23576 18760 23576 18760 0 spi.dout\[6\]
rlabel metal2 26096 19320 26096 19320 0 spi.dout\[7\]
rlabel metal3 37408 23016 37408 23016 0 uart.busy
rlabel metal2 4648 16240 4648 16240 0 uart.counter\[0\]
rlabel metal2 4984 13496 4984 13496 0 uart.counter\[1\]
rlabel metal2 4872 13384 4872 13384 0 uart.counter\[2\]
rlabel metal2 4984 11200 4984 11200 0 uart.counter\[3\]
rlabel metal2 7056 8904 7056 8904 0 uart.data_buff\[0\]
rlabel metal2 9240 11704 9240 11704 0 uart.data_buff\[1\]
rlabel metal2 12992 8904 12992 8904 0 uart.data_buff\[2\]
rlabel metal2 14280 6552 14280 6552 0 uart.data_buff\[3\]
rlabel metal2 16520 9296 16520 9296 0 uart.data_buff\[4\]
rlabel metal2 19880 11760 19880 11760 0 uart.data_buff\[5\]
rlabel metal2 20776 16072 20776 16072 0 uart.data_buff\[6\]
rlabel metal2 18592 18536 18592 18536 0 uart.data_buff\[7\]
rlabel metal2 14728 17920 14728 17920 0 uart.data_buff\[8\]
rlabel metal3 12152 16072 12152 16072 0 uart.data_buff\[9\]
rlabel metal2 8008 25592 8008 25592 0 uart.div_counter\[0\]
rlabel metal2 15176 38080 15176 38080 0 uart.div_counter\[10\]
rlabel metal2 16296 36344 16296 36344 0 uart.div_counter\[11\]
rlabel metal2 14168 30912 14168 30912 0 uart.div_counter\[12\]
rlabel metal2 17752 29792 17752 29792 0 uart.div_counter\[13\]
rlabel metal2 14784 27720 14784 27720 0 uart.div_counter\[14\]
rlabel metal2 14224 24584 14224 24584 0 uart.div_counter\[15\]
rlabel metal2 18872 33096 18872 33096 0 uart.div_counter\[1\]
rlabel metal3 16912 23912 16912 23912 0 uart.div_counter\[2\]
rlabel metal2 16912 32424 16912 32424 0 uart.div_counter\[3\]
rlabel metal2 6440 27496 6440 27496 0 uart.div_counter\[4\]
rlabel metal2 16856 28952 16856 28952 0 uart.div_counter\[5\]
rlabel metal2 15624 30856 15624 30856 0 uart.div_counter\[6\]
rlabel metal3 11088 29624 11088 29624 0 uart.div_counter\[7\]
rlabel metal2 9576 34832 9576 34832 0 uart.div_counter\[8\]
rlabel metal2 18536 35056 18536 35056 0 uart.div_counter\[9\]
rlabel metal2 33320 40320 33320 40320 0 uart.divisor\[0\]
rlabel metal2 24696 36288 24696 36288 0 uart.divisor\[10\]
rlabel metal3 23688 33992 23688 33992 0 uart.divisor\[11\]
rlabel metal2 18200 33656 18200 33656 0 uart.divisor\[12\]
rlabel metal1 17472 38696 17472 38696 0 uart.divisor\[13\]
rlabel metal2 17752 24808 17752 24808 0 uart.divisor\[14\]
rlabel metal2 16744 24808 16744 24808 0 uart.divisor\[15\]
rlabel metal2 21112 38668 21112 38668 0 uart.divisor\[1\]
rlabel metal2 18424 24472 18424 24472 0 uart.divisor\[2\]
rlabel metal2 18424 33376 18424 33376 0 uart.divisor\[3\]
rlabel metal2 17192 27496 17192 27496 0 uart.divisor\[4\]
rlabel metal3 17584 28616 17584 28616 0 uart.divisor\[5\]
rlabel metal2 34440 26656 34440 26656 0 uart.divisor\[6\]
rlabel metal3 29904 26376 29904 26376 0 uart.divisor\[7\]
rlabel metal2 25704 32704 25704 32704 0 uart.divisor\[8\]
rlabel metal2 24696 34608 24696 34608 0 uart.divisor\[9\]
rlabel metal2 38808 37072 38808 37072 0 uart.dout\[0\]
rlabel metal2 39200 34888 39200 34888 0 uart.dout\[1\]
rlabel metal2 36400 39368 36400 39368 0 uart.dout\[2\]
rlabel metal2 44072 41216 44072 41216 0 uart.dout\[3\]
rlabel metal2 44072 38920 44072 38920 0 uart.dout\[4\]
rlabel metal2 46200 39312 46200 39312 0 uart.dout\[5\]
rlabel metal2 42392 36456 42392 36456 0 uart.dout\[6\]
rlabel metal2 40040 40600 40040 40600 0 uart.dout\[7\]
rlabel metal2 41048 26152 41048 26152 0 uart.has_byte
rlabel metal2 39032 46256 39032 46256 0 uart.receive_buff\[0\]
rlabel metal3 37632 48888 37632 48888 0 uart.receive_buff\[1\]
rlabel metal2 41216 50680 41216 50680 0 uart.receive_buff\[2\]
rlabel metal2 45752 47376 45752 47376 0 uart.receive_buff\[3\]
rlabel metal2 44408 44464 44408 44464 0 uart.receive_buff\[4\]
rlabel metal2 43400 45584 43400 45584 0 uart.receive_buff\[5\]
rlabel metal2 43232 42840 43232 42840 0 uart.receive_buff\[6\]
rlabel metal3 40488 45080 40488 45080 0 uart.receive_buff\[7\]
rlabel metal2 48384 50680 48384 50680 0 uart.receive_counter\[0\]
rlabel metal2 53256 46704 53256 46704 0 uart.receive_counter\[1\]
rlabel metal2 53256 49392 53256 49392 0 uart.receive_counter\[2\]
rlabel metal2 49224 44240 49224 44240 0 uart.receive_counter\[3\]
rlabel metal2 24136 42392 24136 42392 0 uart.receive_div_counter\[0\]
rlabel metal4 19096 41216 19096 41216 0 uart.receive_div_counter\[10\]
rlabel metal2 19376 44408 19376 44408 0 uart.receive_div_counter\[11\]
rlabel metal2 12264 44464 12264 44464 0 uart.receive_div_counter\[12\]
rlabel metal2 16968 42560 16968 42560 0 uart.receive_div_counter\[13\]
rlabel metal2 15288 38752 15288 38752 0 uart.receive_div_counter\[14\]
rlabel metal3 15960 39704 15960 39704 0 uart.receive_div_counter\[15\]
rlabel metal2 22512 41160 22512 41160 0 uart.receive_div_counter\[1\]
rlabel metal2 28728 39928 28728 39928 0 uart.receive_div_counter\[2\]
rlabel metal2 24584 41440 24584 41440 0 uart.receive_div_counter\[3\]
rlabel metal2 25032 50428 25032 50428 0 uart.receive_div_counter\[4\]
rlabel metal2 31136 50680 31136 50680 0 uart.receive_div_counter\[5\]
rlabel metal2 30968 46088 30968 46088 0 uart.receive_div_counter\[6\]
rlabel metal2 30296 46704 30296 46704 0 uart.receive_div_counter\[7\]
rlabel metal2 33712 46648 33712 46648 0 uart.receive_div_counter\[8\]
rlabel metal2 18592 50680 18592 50680 0 uart.receive_div_counter\[9\]
rlabel metal2 35560 45080 35560 45080 0 uart.receiving
rlabel metal2 39592 29568 39592 29568 0 uart_ien
rlabel metal2 22792 47096 22792 47096 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 55000 55000
<< end >>
